magic
tech sky130A
magscale 1 2
timestamp 1725110490
<< viali >>
rect 1397 6772 1431 11864
rect 2769 6772 2803 11864
<< metal1 >>
rect 4188 33680 4246 33686
rect 4188 33628 4191 33680
rect 4243 33628 4246 33680
rect 4188 33600 4246 33628
rect 4194 33246 4240 33600
rect 4076 33200 4240 33246
rect 3932 32934 3990 33084
rect 3340 32168 3610 32218
rect 3340 31680 3390 32168
rect 4194 32010 4240 33200
rect 4086 31964 4240 32010
rect 4073 31391 4125 31397
rect 561 31253 619 31259
rect 561 31201 564 31253
rect 616 31201 619 31253
rect 561 31052 619 31201
rect 189 30839 241 30845
rect 189 19465 241 19471
rect 4073 19021 4125 19027
rect 1391 12036 1484 12082
rect 2716 12036 2809 12082
rect 1391 11864 1437 12036
rect 1391 6772 1397 11864
rect 1431 6772 1437 11864
rect 1576 11722 1669 12035
rect 2531 11722 2624 12035
rect 2763 11864 2809 12036
rect 1391 6760 1437 6772
rect 2763 6772 2769 11864
rect 2803 6772 2809 11864
rect 2763 6760 2809 6772
<< via1 >>
rect 4191 33628 4243 33680
rect 4030 33302 4150 33474
rect 4030 33090 4150 33146
rect 3764 32826 3960 32894
rect 3458 32384 3808 32560
rect 3764 32050 3960 32118
rect 564 31201 616 31253
rect 189 19471 241 30839
rect 4073 19027 4125 31391
rect 1537 6914 2663 7323
<< metal2 >>
rect 4189 33682 4245 33691
rect 4189 33617 4245 33626
rect 4030 33474 4150 33480
rect 4030 33296 4150 33302
rect 3898 33146 4150 33152
rect 3898 33143 4030 33146
rect 3898 32894 3903 33143
rect 3961 33090 4030 33143
rect 3961 33084 4150 33090
rect 3758 32826 3764 32894
rect 3452 32384 3458 32560
rect 3808 32384 3814 32560
rect 3898 32118 3903 32826
rect 3758 32050 3764 32118
rect 3961 32059 3966 33084
rect 3960 32050 3966 32059
rect 3240 31546 3297 31555
rect 562 31255 618 31264
rect 562 31190 618 31199
rect 189 30839 381 30845
rect 241 19471 381 30839
rect 189 19465 381 19471
rect 3897 31391 4125 31397
rect 3897 19027 4073 31391
rect 3897 19021 4125 19027
rect 3240 18863 3297 18872
rect 1531 6914 1537 7323
rect 2663 6914 2669 7323
<< via2 >>
rect 4189 33680 4245 33682
rect 4189 33628 4191 33680
rect 4191 33628 4243 33680
rect 4243 33628 4245 33680
rect 4189 33626 4245 33628
rect 4035 33305 4093 33471
rect 3903 32894 3961 33143
rect 3903 32826 3960 32894
rect 3960 32826 3961 32894
rect 3461 32389 3805 32555
rect 3903 32118 3961 32826
rect 3903 32059 3960 32118
rect 3960 32059 3961 32118
rect 562 31253 618 31255
rect 562 31201 564 31253
rect 564 31201 616 31253
rect 616 31201 618 31253
rect 562 31199 618 31201
rect 386 19474 616 30836
rect 746 19378 981 30932
rect 3240 18872 3532 31546
rect 3662 19030 3892 31388
rect 1540 6919 2660 7318
<< metal3 >>
rect 1000 38499 4098 38500
rect 1000 38433 1006 38499
rect 1599 38433 4098 38499
rect 1000 38432 4098 38433
rect 1800 38359 3966 38360
rect 1800 38293 1806 38359
rect 2399 38293 3966 38359
rect 1800 38292 3966 38293
rect 962 31300 1400 38144
rect 542 31259 638 31277
rect 542 31195 558 31259
rect 622 31195 638 31259
rect 542 31177 638 31195
rect 960 30941 1400 31300
rect 741 30932 1400 30941
rect 381 30839 621 30845
rect 381 19471 382 30839
rect 620 19471 621 30839
rect 381 19465 621 19471
rect 741 19378 746 30932
rect 981 19378 1400 30932
rect 741 19369 1400 19378
rect 960 12166 1400 19369
rect 2800 31580 3240 38144
rect 3898 33143 3966 38292
rect 4030 33471 4098 38432
rect 4169 33686 4265 33704
rect 4169 33622 4185 33686
rect 4249 33622 4265 33686
rect 4169 33604 4265 33622
rect 4030 33305 4035 33471
rect 4093 33305 4098 33471
rect 4030 33296 4098 33305
rect 3452 32559 3814 32560
rect 3452 32385 3458 32559
rect 3808 32385 3814 32559
rect 3452 32384 3814 32385
rect 3898 32059 3903 33143
rect 3961 32059 3966 33143
rect 3898 32050 3966 32059
rect 2800 31546 3537 31580
rect 2800 18872 3240 31546
rect 3532 18872 3537 31546
rect 3657 31391 3897 31397
rect 3657 19027 3658 31391
rect 3896 19027 3897 31391
rect 3657 19021 3897 19027
rect 2800 18840 3537 18872
rect 2800 12166 3240 18840
rect 1531 7318 2669 7323
rect 1531 6919 1540 7318
rect 2660 6919 2669 7318
rect 1531 6914 2669 6919
rect 2489 2180 2669 6914
rect 2489 2179 3800 2180
rect 2489 2001 3446 2179
rect 3614 2178 3800 2179
rect 3794 2001 3800 2178
rect 2489 2000 3800 2001
<< via3 >>
rect 1006 38433 1599 38499
rect 1806 38293 2399 38359
rect 558 31255 622 31259
rect 558 31199 562 31255
rect 562 31199 618 31255
rect 618 31199 622 31255
rect 558 31195 622 31199
rect 382 30836 620 30839
rect 382 19474 386 30836
rect 386 19474 616 30836
rect 616 19474 620 30836
rect 382 19471 620 19474
rect 1801 12172 2399 38138
rect 4185 33682 4249 33686
rect 4185 33626 4189 33682
rect 4189 33626 4245 33682
rect 4245 33626 4249 33682
rect 4185 33622 4249 33626
rect 3458 32555 3808 32559
rect 3458 32389 3461 32555
rect 3461 32389 3805 32555
rect 3805 32389 3808 32555
rect 3458 32385 3808 32389
rect 3658 31388 3896 31391
rect 3658 19030 3662 31388
rect 3662 19030 3892 31388
rect 3892 19030 3896 31388
rect 3658 19027 3896 19030
rect 3446 2178 3614 2179
rect 3446 2001 3794 2178
<< metal4 >>
rect 3006 44952 3066 45152
rect 3558 44952 3618 45152
rect 4110 44952 4170 45152
rect 4662 44952 4722 45152
rect 5214 44952 5274 45152
rect 5766 44952 5826 45152
rect 6318 44952 6378 45152
rect 6870 44952 6930 45152
rect 3006 44892 6930 44952
rect 7422 44952 7482 45152
rect 7974 44952 8034 45152
rect 8526 44952 8586 45152
rect 9078 44952 9138 45152
rect 9630 44952 9690 45152
rect 10182 44952 10242 45152
rect 10734 44952 10794 45152
rect 11286 44952 11346 45152
rect 11838 44952 11898 45152
rect 12390 44952 12450 45152
rect 12942 44952 13002 45152
rect 13494 44952 13554 45152
rect 14046 44952 14106 45152
rect 14598 44952 14658 45152
rect 15150 44952 15210 45152
rect 15702 44952 15762 45152
rect 16254 44952 16314 45152
rect 16806 44952 16866 45152
rect 17358 44952 17418 45152
rect 17910 44952 17970 45152
rect 18462 44952 18522 45152
rect 19014 44952 19074 45152
rect 19566 44952 19626 45152
rect 20118 44952 20178 45152
rect 7422 44892 15762 44952
rect 6870 44720 6930 44892
rect 15702 44860 15762 44892
rect 20670 44860 20730 45152
rect 15702 44800 20730 44860
rect 21222 44720 21282 45152
rect 21774 44952 21834 45152
rect 22326 44952 22386 45152
rect 22878 44952 22938 45152
rect 23430 44952 23490 45152
rect 6870 44660 21282 44720
rect 23982 44580 24042 45152
rect 560 44520 24042 44580
rect 560 31260 620 44520
rect 24534 44440 24594 45152
rect 25086 44952 25146 45152
rect 25638 44952 25698 45152
rect 26190 44952 26250 45152
rect 4187 44380 24594 44440
rect 1000 38499 1600 44152
rect 1000 38433 1006 38499
rect 1599 38433 1600 38499
rect 557 31259 623 31260
rect 557 31195 558 31259
rect 622 31195 623 31259
rect 557 31194 623 31195
rect 1000 30845 1600 38433
rect 381 30839 1600 30845
rect 381 19471 382 30839
rect 620 19471 1600 30839
rect 381 19465 1600 19471
rect 1000 980 1600 19465
rect 1800 38359 2400 44152
rect 1800 38293 1806 38359
rect 2399 38293 2400 38359
rect 1800 38138 2400 38293
rect 1800 12172 1801 38138
rect 2399 12172 2400 38138
rect 1800 1380 2400 12172
rect 2600 32560 3200 44152
rect 4187 33687 4247 44380
rect 4184 33686 4250 33687
rect 4184 33622 4185 33686
rect 4249 33622 4250 33686
rect 4184 33621 4250 33622
rect 2600 32559 3814 32560
rect 2600 32385 3458 32559
rect 3808 32385 3814 32559
rect 2600 32384 3814 32385
rect 2600 31397 3200 32384
rect 2600 31391 3897 31397
rect 2600 19027 3658 31391
rect 3896 19027 3897 31391
rect 2600 19021 3897 19027
rect 2600 1780 3200 19021
rect 3440 2179 27414 2180
rect 3440 2001 3446 2179
rect 3614 2178 27414 2179
rect 3794 2001 27414 2178
rect 3440 2000 27414 2001
rect 2600 1600 23550 1780
rect 1798 1200 19686 1380
rect 1000 800 15822 980
rect 7914 300 11958 480
rect 186 0 366 200
rect 4050 0 4230 200
rect 7914 0 8094 300
rect 11778 0 11958 300
rect 15642 0 15822 800
rect 19506 0 19686 1200
rect 23370 0 23550 1600
rect 27234 0 27414 2000
use inv  inv_0
timestamp 1725098041
transform -1 0 4840 0 -1 38368
box 668 4844 940 5328
use lv2hv  lv2hv_0
timestamp 1725098041
transform 1 0 3382 0 1 32472
box -2 -532 804 532
use nfet_load  nfet_load_0
timestamp 1725098041
transform 0 1 2100 -1 0 25155
box -13155 -700 13155 700
use pfet_vapwr  pfet_vapwr_0
timestamp 1725098041
transform 0 1 3597 -1 0 25209
box -6549 -597 6549 597
use pfet_vdpwr  pfet_vdpwr_0
timestamp 1725098041
transform 0 -1 681 -1 0 25155
box -5927 -519 5927 519
use res_bias  res_bias_0
timestamp 1725098041
transform -1 0 2100 0 -1 9318
box -739 -2582 739 2582
<< labels >>
flabel metal4 s 25638 44952 25698 45152 0 FreeSans 480 90 0 0 clk
port 0 nsew signal input
flabel metal4 s 26190 44952 26250 45152 0 FreeSans 480 90 0 0 ena
port 1 nsew signal input
flabel metal4 s 25086 44952 25146 45152 0 FreeSans 480 90 0 0 rst_n
port 2 nsew signal input
flabel metal4 s 27234 0 27414 200 0 FreeSans 960 0 0 0 ua[0]
port 3 nsew signal bidirectional
flabel metal4 s 23370 0 23550 200 0 FreeSans 960 0 0 0 ua[1]
port 4 nsew signal bidirectional
flabel metal4 s 19506 0 19686 200 0 FreeSans 960 0 0 0 ua[2]
port 5 nsew signal bidirectional
flabel metal4 s 15642 0 15822 200 0 FreeSans 960 0 0 0 ua[3]
port 6 nsew signal bidirectional
flabel metal4 s 11778 0 11958 200 0 FreeSans 960 0 0 0 ua[4]
port 7 nsew signal bidirectional
flabel metal4 s 7914 0 8094 200 0 FreeSans 960 0 0 0 ua[5]
port 8 nsew signal bidirectional
flabel metal4 s 4050 0 4230 200 0 FreeSans 960 0 0 0 ua[6]
port 9 nsew signal bidirectional
flabel metal4 s 186 0 366 200 0 FreeSans 960 0 0 0 ua[7]
port 10 nsew signal bidirectional
flabel metal4 s 24534 44952 24594 45152 0 FreeSans 480 90 0 0 ui_in[0]
port 11 nsew signal input
flabel metal4 s 23982 44952 24042 45152 0 FreeSans 480 90 0 0 ui_in[1]
port 12 nsew signal input
flabel metal4 s 23430 44952 23490 45152 0 FreeSans 480 90 0 0 ui_in[2]
port 13 nsew signal input
flabel metal4 s 22878 44952 22938 45152 0 FreeSans 480 90 0 0 ui_in[3]
port 14 nsew signal input
flabel metal4 s 22326 44952 22386 45152 0 FreeSans 480 90 0 0 ui_in[4]
port 15 nsew signal input
flabel metal4 s 21774 44952 21834 45152 0 FreeSans 480 90 0 0 ui_in[5]
port 16 nsew signal input
flabel metal4 s 21222 44952 21282 45152 0 FreeSans 480 90 0 0 ui_in[6]
port 17 nsew signal input
flabel metal4 s 20670 44952 20730 45152 0 FreeSans 480 90 0 0 ui_in[7]
port 18 nsew signal input
flabel metal4 s 20118 44952 20178 45152 0 FreeSans 480 90 0 0 uio_in[0]
port 19 nsew signal input
flabel metal4 s 19566 44952 19626 45152 0 FreeSans 480 90 0 0 uio_in[1]
port 20 nsew signal input
flabel metal4 s 19014 44952 19074 45152 0 FreeSans 480 90 0 0 uio_in[2]
port 21 nsew signal input
flabel metal4 s 18462 44952 18522 45152 0 FreeSans 480 90 0 0 uio_in[3]
port 22 nsew signal input
flabel metal4 s 17910 44952 17970 45152 0 FreeSans 480 90 0 0 uio_in[4]
port 23 nsew signal input
flabel metal4 s 17358 44952 17418 45152 0 FreeSans 480 90 0 0 uio_in[5]
port 24 nsew signal input
flabel metal4 s 16806 44952 16866 45152 0 FreeSans 480 90 0 0 uio_in[6]
port 25 nsew signal input
flabel metal4 s 16254 44952 16314 45152 0 FreeSans 480 90 0 0 uio_in[7]
port 26 nsew signal input
flabel metal4 s 6870 44952 6930 45152 0 FreeSans 480 90 0 0 uio_oe[0]
port 27 nsew signal output
flabel metal4 s 6318 44952 6378 45152 0 FreeSans 480 90 0 0 uio_oe[1]
port 28 nsew signal output
flabel metal4 s 5766 44952 5826 45152 0 FreeSans 480 90 0 0 uio_oe[2]
port 29 nsew signal output
flabel metal4 s 5214 44952 5274 45152 0 FreeSans 480 90 0 0 uio_oe[3]
port 30 nsew signal output
flabel metal4 s 4662 44952 4722 45152 0 FreeSans 480 90 0 0 uio_oe[4]
port 31 nsew signal output
flabel metal4 s 4110 44952 4170 45152 0 FreeSans 480 90 0 0 uio_oe[5]
port 32 nsew signal output
flabel metal4 s 3558 44952 3618 45152 0 FreeSans 480 90 0 0 uio_oe[6]
port 33 nsew signal output
flabel metal4 s 3006 44952 3066 45152 0 FreeSans 480 90 0 0 uio_oe[7]
port 34 nsew signal output
flabel metal4 s 11286 44952 11346 45152 0 FreeSans 480 90 0 0 uio_out[0]
port 35 nsew signal output
flabel metal4 s 10734 44952 10794 45152 0 FreeSans 480 90 0 0 uio_out[1]
port 36 nsew signal output
flabel metal4 s 10182 44952 10242 45152 0 FreeSans 480 90 0 0 uio_out[2]
port 37 nsew signal output
flabel metal4 s 9630 44952 9690 45152 0 FreeSans 480 90 0 0 uio_out[3]
port 38 nsew signal output
flabel metal4 s 9078 44952 9138 45152 0 FreeSans 480 90 0 0 uio_out[4]
port 39 nsew signal output
flabel metal4 s 8526 44952 8586 45152 0 FreeSans 480 90 0 0 uio_out[5]
port 40 nsew signal output
flabel metal4 s 7974 44952 8034 45152 0 FreeSans 480 90 0 0 uio_out[6]
port 41 nsew signal output
flabel metal4 s 7422 44952 7482 45152 0 FreeSans 480 90 0 0 uio_out[7]
port 42 nsew signal output
flabel metal4 s 15702 44952 15762 45152 0 FreeSans 480 90 0 0 uo_out[0]
port 43 nsew signal output
flabel metal4 s 15150 44952 15210 45152 0 FreeSans 480 90 0 0 uo_out[1]
port 44 nsew signal output
flabel metal4 s 14598 44952 14658 45152 0 FreeSans 480 90 0 0 uo_out[2]
port 45 nsew signal output
flabel metal4 s 14046 44952 14106 45152 0 FreeSans 480 90 0 0 uo_out[3]
port 46 nsew signal output
flabel metal4 s 13494 44952 13554 45152 0 FreeSans 480 90 0 0 uo_out[4]
port 47 nsew signal output
flabel metal4 s 12942 44952 13002 45152 0 FreeSans 480 90 0 0 uo_out[5]
port 48 nsew signal output
flabel metal4 s 12390 44952 12450 45152 0 FreeSans 480 90 0 0 uo_out[6]
port 49 nsew signal output
flabel metal4 s 11838 44952 11898 45152 0 FreeSans 480 90 0 0 uo_out[7]
port 50 nsew signal output
flabel metal4 s 1800 1200 2400 44152 0 FreeSans 160 0 0 0 VGND
port 51 nsew
flabel metal4 s 1000 800 1600 44152 0 FreeSans 160 0 0 0 VDPWR
port 52 nsew
flabel metal4 s 2600 1600 3200 44152 0 FreeSans 160 0 0 0 VAPWR
port 53 nsew
<< properties >>
string FIXED_BBOX 0 0 29072 45152
<< end >>
