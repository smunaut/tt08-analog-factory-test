magic
tech sky130A
magscale 1 2
timestamp 1725098041
<< nwell >>
rect -5927 -519 5927 519
<< pmos >>
rect -5727 -300 -5697 300
rect -5631 -300 -5601 300
rect -5535 -300 -5505 300
rect -5439 -300 -5409 300
rect -5343 -300 -5313 300
rect -5247 -300 -5217 300
rect -5151 -300 -5121 300
rect -5055 -300 -5025 300
rect -4959 -300 -4929 300
rect -4863 -300 -4833 300
rect -4767 -300 -4737 300
rect -4671 -300 -4641 300
rect -4575 -300 -4545 300
rect -4479 -300 -4449 300
rect -4383 -300 -4353 300
rect -4287 -300 -4257 300
rect -4191 -300 -4161 300
rect -4095 -300 -4065 300
rect -3999 -300 -3969 300
rect -3903 -300 -3873 300
rect -3807 -300 -3777 300
rect -3711 -300 -3681 300
rect -3615 -300 -3585 300
rect -3519 -300 -3489 300
rect -3423 -300 -3393 300
rect -3327 -300 -3297 300
rect -3231 -300 -3201 300
rect -3135 -300 -3105 300
rect -3039 -300 -3009 300
rect -2943 -300 -2913 300
rect -2847 -300 -2817 300
rect -2751 -300 -2721 300
rect -2655 -300 -2625 300
rect -2559 -300 -2529 300
rect -2463 -300 -2433 300
rect -2367 -300 -2337 300
rect -2271 -300 -2241 300
rect -2175 -300 -2145 300
rect -2079 -300 -2049 300
rect -1983 -300 -1953 300
rect -1887 -300 -1857 300
rect -1791 -300 -1761 300
rect -1695 -300 -1665 300
rect -1599 -300 -1569 300
rect -1503 -300 -1473 300
rect -1407 -300 -1377 300
rect -1311 -300 -1281 300
rect -1215 -300 -1185 300
rect -1119 -300 -1089 300
rect -1023 -300 -993 300
rect -927 -300 -897 300
rect -831 -300 -801 300
rect -735 -300 -705 300
rect -639 -300 -609 300
rect -543 -300 -513 300
rect -447 -300 -417 300
rect -351 -300 -321 300
rect -255 -300 -225 300
rect -159 -300 -129 300
rect -63 -300 -33 300
rect 33 -300 63 300
rect 129 -300 159 300
rect 225 -300 255 300
rect 321 -300 351 300
rect 417 -300 447 300
rect 513 -300 543 300
rect 609 -300 639 300
rect 705 -300 735 300
rect 801 -300 831 300
rect 897 -300 927 300
rect 993 -300 1023 300
rect 1089 -300 1119 300
rect 1185 -300 1215 300
rect 1281 -300 1311 300
rect 1377 -300 1407 300
rect 1473 -300 1503 300
rect 1569 -300 1599 300
rect 1665 -300 1695 300
rect 1761 -300 1791 300
rect 1857 -300 1887 300
rect 1953 -300 1983 300
rect 2049 -300 2079 300
rect 2145 -300 2175 300
rect 2241 -300 2271 300
rect 2337 -300 2367 300
rect 2433 -300 2463 300
rect 2529 -300 2559 300
rect 2625 -300 2655 300
rect 2721 -300 2751 300
rect 2817 -300 2847 300
rect 2913 -300 2943 300
rect 3009 -300 3039 300
rect 3105 -300 3135 300
rect 3201 -300 3231 300
rect 3297 -300 3327 300
rect 3393 -300 3423 300
rect 3489 -300 3519 300
rect 3585 -300 3615 300
rect 3681 -300 3711 300
rect 3777 -300 3807 300
rect 3873 -300 3903 300
rect 3969 -300 3999 300
rect 4065 -300 4095 300
rect 4161 -300 4191 300
rect 4257 -300 4287 300
rect 4353 -300 4383 300
rect 4449 -300 4479 300
rect 4545 -300 4575 300
rect 4641 -300 4671 300
rect 4737 -300 4767 300
rect 4833 -300 4863 300
rect 4929 -300 4959 300
rect 5025 -300 5055 300
rect 5121 -300 5151 300
rect 5217 -300 5247 300
rect 5313 -300 5343 300
rect 5409 -300 5439 300
rect 5505 -300 5535 300
rect 5601 -300 5631 300
rect 5697 -300 5727 300
<< pdiff >>
rect -5789 288 -5727 300
rect -5789 -288 -5777 288
rect -5743 -288 -5727 288
rect -5789 -300 -5727 -288
rect -5697 288 -5631 300
rect -5697 -288 -5681 288
rect -5647 -288 -5631 288
rect -5697 -300 -5631 -288
rect -5601 288 -5535 300
rect -5601 -288 -5585 288
rect -5551 -288 -5535 288
rect -5601 -300 -5535 -288
rect -5505 288 -5439 300
rect -5505 -288 -5489 288
rect -5455 -288 -5439 288
rect -5505 -300 -5439 -288
rect -5409 288 -5343 300
rect -5409 -288 -5393 288
rect -5359 -288 -5343 288
rect -5409 -300 -5343 -288
rect -5313 288 -5247 300
rect -5313 -288 -5297 288
rect -5263 -288 -5247 288
rect -5313 -300 -5247 -288
rect -5217 288 -5151 300
rect -5217 -288 -5201 288
rect -5167 -288 -5151 288
rect -5217 -300 -5151 -288
rect -5121 288 -5055 300
rect -5121 -288 -5105 288
rect -5071 -288 -5055 288
rect -5121 -300 -5055 -288
rect -5025 288 -4959 300
rect -5025 -288 -5009 288
rect -4975 -288 -4959 288
rect -5025 -300 -4959 -288
rect -4929 288 -4863 300
rect -4929 -288 -4913 288
rect -4879 -288 -4863 288
rect -4929 -300 -4863 -288
rect -4833 288 -4767 300
rect -4833 -288 -4817 288
rect -4783 -288 -4767 288
rect -4833 -300 -4767 -288
rect -4737 288 -4671 300
rect -4737 -288 -4721 288
rect -4687 -288 -4671 288
rect -4737 -300 -4671 -288
rect -4641 288 -4575 300
rect -4641 -288 -4625 288
rect -4591 -288 -4575 288
rect -4641 -300 -4575 -288
rect -4545 288 -4479 300
rect -4545 -288 -4529 288
rect -4495 -288 -4479 288
rect -4545 -300 -4479 -288
rect -4449 288 -4383 300
rect -4449 -288 -4433 288
rect -4399 -288 -4383 288
rect -4449 -300 -4383 -288
rect -4353 288 -4287 300
rect -4353 -288 -4337 288
rect -4303 -288 -4287 288
rect -4353 -300 -4287 -288
rect -4257 288 -4191 300
rect -4257 -288 -4241 288
rect -4207 -288 -4191 288
rect -4257 -300 -4191 -288
rect -4161 288 -4095 300
rect -4161 -288 -4145 288
rect -4111 -288 -4095 288
rect -4161 -300 -4095 -288
rect -4065 288 -3999 300
rect -4065 -288 -4049 288
rect -4015 -288 -3999 288
rect -4065 -300 -3999 -288
rect -3969 288 -3903 300
rect -3969 -288 -3953 288
rect -3919 -288 -3903 288
rect -3969 -300 -3903 -288
rect -3873 288 -3807 300
rect -3873 -288 -3857 288
rect -3823 -288 -3807 288
rect -3873 -300 -3807 -288
rect -3777 288 -3711 300
rect -3777 -288 -3761 288
rect -3727 -288 -3711 288
rect -3777 -300 -3711 -288
rect -3681 288 -3615 300
rect -3681 -288 -3665 288
rect -3631 -288 -3615 288
rect -3681 -300 -3615 -288
rect -3585 288 -3519 300
rect -3585 -288 -3569 288
rect -3535 -288 -3519 288
rect -3585 -300 -3519 -288
rect -3489 288 -3423 300
rect -3489 -288 -3473 288
rect -3439 -288 -3423 288
rect -3489 -300 -3423 -288
rect -3393 288 -3327 300
rect -3393 -288 -3377 288
rect -3343 -288 -3327 288
rect -3393 -300 -3327 -288
rect -3297 288 -3231 300
rect -3297 -288 -3281 288
rect -3247 -288 -3231 288
rect -3297 -300 -3231 -288
rect -3201 288 -3135 300
rect -3201 -288 -3185 288
rect -3151 -288 -3135 288
rect -3201 -300 -3135 -288
rect -3105 288 -3039 300
rect -3105 -288 -3089 288
rect -3055 -288 -3039 288
rect -3105 -300 -3039 -288
rect -3009 288 -2943 300
rect -3009 -288 -2993 288
rect -2959 -288 -2943 288
rect -3009 -300 -2943 -288
rect -2913 288 -2847 300
rect -2913 -288 -2897 288
rect -2863 -288 -2847 288
rect -2913 -300 -2847 -288
rect -2817 288 -2751 300
rect -2817 -288 -2801 288
rect -2767 -288 -2751 288
rect -2817 -300 -2751 -288
rect -2721 288 -2655 300
rect -2721 -288 -2705 288
rect -2671 -288 -2655 288
rect -2721 -300 -2655 -288
rect -2625 288 -2559 300
rect -2625 -288 -2609 288
rect -2575 -288 -2559 288
rect -2625 -300 -2559 -288
rect -2529 288 -2463 300
rect -2529 -288 -2513 288
rect -2479 -288 -2463 288
rect -2529 -300 -2463 -288
rect -2433 288 -2367 300
rect -2433 -288 -2417 288
rect -2383 -288 -2367 288
rect -2433 -300 -2367 -288
rect -2337 288 -2271 300
rect -2337 -288 -2321 288
rect -2287 -288 -2271 288
rect -2337 -300 -2271 -288
rect -2241 288 -2175 300
rect -2241 -288 -2225 288
rect -2191 -288 -2175 288
rect -2241 -300 -2175 -288
rect -2145 288 -2079 300
rect -2145 -288 -2129 288
rect -2095 -288 -2079 288
rect -2145 -300 -2079 -288
rect -2049 288 -1983 300
rect -2049 -288 -2033 288
rect -1999 -288 -1983 288
rect -2049 -300 -1983 -288
rect -1953 288 -1887 300
rect -1953 -288 -1937 288
rect -1903 -288 -1887 288
rect -1953 -300 -1887 -288
rect -1857 288 -1791 300
rect -1857 -288 -1841 288
rect -1807 -288 -1791 288
rect -1857 -300 -1791 -288
rect -1761 288 -1695 300
rect -1761 -288 -1745 288
rect -1711 -288 -1695 288
rect -1761 -300 -1695 -288
rect -1665 288 -1599 300
rect -1665 -288 -1649 288
rect -1615 -288 -1599 288
rect -1665 -300 -1599 -288
rect -1569 288 -1503 300
rect -1569 -288 -1553 288
rect -1519 -288 -1503 288
rect -1569 -300 -1503 -288
rect -1473 288 -1407 300
rect -1473 -288 -1457 288
rect -1423 -288 -1407 288
rect -1473 -300 -1407 -288
rect -1377 288 -1311 300
rect -1377 -288 -1361 288
rect -1327 -288 -1311 288
rect -1377 -300 -1311 -288
rect -1281 288 -1215 300
rect -1281 -288 -1265 288
rect -1231 -288 -1215 288
rect -1281 -300 -1215 -288
rect -1185 288 -1119 300
rect -1185 -288 -1169 288
rect -1135 -288 -1119 288
rect -1185 -300 -1119 -288
rect -1089 288 -1023 300
rect -1089 -288 -1073 288
rect -1039 -288 -1023 288
rect -1089 -300 -1023 -288
rect -993 288 -927 300
rect -993 -288 -977 288
rect -943 -288 -927 288
rect -993 -300 -927 -288
rect -897 288 -831 300
rect -897 -288 -881 288
rect -847 -288 -831 288
rect -897 -300 -831 -288
rect -801 288 -735 300
rect -801 -288 -785 288
rect -751 -288 -735 288
rect -801 -300 -735 -288
rect -705 288 -639 300
rect -705 -288 -689 288
rect -655 -288 -639 288
rect -705 -300 -639 -288
rect -609 288 -543 300
rect -609 -288 -593 288
rect -559 -288 -543 288
rect -609 -300 -543 -288
rect -513 288 -447 300
rect -513 -288 -497 288
rect -463 -288 -447 288
rect -513 -300 -447 -288
rect -417 288 -351 300
rect -417 -288 -401 288
rect -367 -288 -351 288
rect -417 -300 -351 -288
rect -321 288 -255 300
rect -321 -288 -305 288
rect -271 -288 -255 288
rect -321 -300 -255 -288
rect -225 288 -159 300
rect -225 -288 -209 288
rect -175 -288 -159 288
rect -225 -300 -159 -288
rect -129 288 -63 300
rect -129 -288 -113 288
rect -79 -288 -63 288
rect -129 -300 -63 -288
rect -33 288 33 300
rect -33 -288 -17 288
rect 17 -288 33 288
rect -33 -300 33 -288
rect 63 288 129 300
rect 63 -288 79 288
rect 113 -288 129 288
rect 63 -300 129 -288
rect 159 288 225 300
rect 159 -288 175 288
rect 209 -288 225 288
rect 159 -300 225 -288
rect 255 288 321 300
rect 255 -288 271 288
rect 305 -288 321 288
rect 255 -300 321 -288
rect 351 288 417 300
rect 351 -288 367 288
rect 401 -288 417 288
rect 351 -300 417 -288
rect 447 288 513 300
rect 447 -288 463 288
rect 497 -288 513 288
rect 447 -300 513 -288
rect 543 288 609 300
rect 543 -288 559 288
rect 593 -288 609 288
rect 543 -300 609 -288
rect 639 288 705 300
rect 639 -288 655 288
rect 689 -288 705 288
rect 639 -300 705 -288
rect 735 288 801 300
rect 735 -288 751 288
rect 785 -288 801 288
rect 735 -300 801 -288
rect 831 288 897 300
rect 831 -288 847 288
rect 881 -288 897 288
rect 831 -300 897 -288
rect 927 288 993 300
rect 927 -288 943 288
rect 977 -288 993 288
rect 927 -300 993 -288
rect 1023 288 1089 300
rect 1023 -288 1039 288
rect 1073 -288 1089 288
rect 1023 -300 1089 -288
rect 1119 288 1185 300
rect 1119 -288 1135 288
rect 1169 -288 1185 288
rect 1119 -300 1185 -288
rect 1215 288 1281 300
rect 1215 -288 1231 288
rect 1265 -288 1281 288
rect 1215 -300 1281 -288
rect 1311 288 1377 300
rect 1311 -288 1327 288
rect 1361 -288 1377 288
rect 1311 -300 1377 -288
rect 1407 288 1473 300
rect 1407 -288 1423 288
rect 1457 -288 1473 288
rect 1407 -300 1473 -288
rect 1503 288 1569 300
rect 1503 -288 1519 288
rect 1553 -288 1569 288
rect 1503 -300 1569 -288
rect 1599 288 1665 300
rect 1599 -288 1615 288
rect 1649 -288 1665 288
rect 1599 -300 1665 -288
rect 1695 288 1761 300
rect 1695 -288 1711 288
rect 1745 -288 1761 288
rect 1695 -300 1761 -288
rect 1791 288 1857 300
rect 1791 -288 1807 288
rect 1841 -288 1857 288
rect 1791 -300 1857 -288
rect 1887 288 1953 300
rect 1887 -288 1903 288
rect 1937 -288 1953 288
rect 1887 -300 1953 -288
rect 1983 288 2049 300
rect 1983 -288 1999 288
rect 2033 -288 2049 288
rect 1983 -300 2049 -288
rect 2079 288 2145 300
rect 2079 -288 2095 288
rect 2129 -288 2145 288
rect 2079 -300 2145 -288
rect 2175 288 2241 300
rect 2175 -288 2191 288
rect 2225 -288 2241 288
rect 2175 -300 2241 -288
rect 2271 288 2337 300
rect 2271 -288 2287 288
rect 2321 -288 2337 288
rect 2271 -300 2337 -288
rect 2367 288 2433 300
rect 2367 -288 2383 288
rect 2417 -288 2433 288
rect 2367 -300 2433 -288
rect 2463 288 2529 300
rect 2463 -288 2479 288
rect 2513 -288 2529 288
rect 2463 -300 2529 -288
rect 2559 288 2625 300
rect 2559 -288 2575 288
rect 2609 -288 2625 288
rect 2559 -300 2625 -288
rect 2655 288 2721 300
rect 2655 -288 2671 288
rect 2705 -288 2721 288
rect 2655 -300 2721 -288
rect 2751 288 2817 300
rect 2751 -288 2767 288
rect 2801 -288 2817 288
rect 2751 -300 2817 -288
rect 2847 288 2913 300
rect 2847 -288 2863 288
rect 2897 -288 2913 288
rect 2847 -300 2913 -288
rect 2943 288 3009 300
rect 2943 -288 2959 288
rect 2993 -288 3009 288
rect 2943 -300 3009 -288
rect 3039 288 3105 300
rect 3039 -288 3055 288
rect 3089 -288 3105 288
rect 3039 -300 3105 -288
rect 3135 288 3201 300
rect 3135 -288 3151 288
rect 3185 -288 3201 288
rect 3135 -300 3201 -288
rect 3231 288 3297 300
rect 3231 -288 3247 288
rect 3281 -288 3297 288
rect 3231 -300 3297 -288
rect 3327 288 3393 300
rect 3327 -288 3343 288
rect 3377 -288 3393 288
rect 3327 -300 3393 -288
rect 3423 288 3489 300
rect 3423 -288 3439 288
rect 3473 -288 3489 288
rect 3423 -300 3489 -288
rect 3519 288 3585 300
rect 3519 -288 3535 288
rect 3569 -288 3585 288
rect 3519 -300 3585 -288
rect 3615 288 3681 300
rect 3615 -288 3631 288
rect 3665 -288 3681 288
rect 3615 -300 3681 -288
rect 3711 288 3777 300
rect 3711 -288 3727 288
rect 3761 -288 3777 288
rect 3711 -300 3777 -288
rect 3807 288 3873 300
rect 3807 -288 3823 288
rect 3857 -288 3873 288
rect 3807 -300 3873 -288
rect 3903 288 3969 300
rect 3903 -288 3919 288
rect 3953 -288 3969 288
rect 3903 -300 3969 -288
rect 3999 288 4065 300
rect 3999 -288 4015 288
rect 4049 -288 4065 288
rect 3999 -300 4065 -288
rect 4095 288 4161 300
rect 4095 -288 4111 288
rect 4145 -288 4161 288
rect 4095 -300 4161 -288
rect 4191 288 4257 300
rect 4191 -288 4207 288
rect 4241 -288 4257 288
rect 4191 -300 4257 -288
rect 4287 288 4353 300
rect 4287 -288 4303 288
rect 4337 -288 4353 288
rect 4287 -300 4353 -288
rect 4383 288 4449 300
rect 4383 -288 4399 288
rect 4433 -288 4449 288
rect 4383 -300 4449 -288
rect 4479 288 4545 300
rect 4479 -288 4495 288
rect 4529 -288 4545 288
rect 4479 -300 4545 -288
rect 4575 288 4641 300
rect 4575 -288 4591 288
rect 4625 -288 4641 288
rect 4575 -300 4641 -288
rect 4671 288 4737 300
rect 4671 -288 4687 288
rect 4721 -288 4737 288
rect 4671 -300 4737 -288
rect 4767 288 4833 300
rect 4767 -288 4783 288
rect 4817 -288 4833 288
rect 4767 -300 4833 -288
rect 4863 288 4929 300
rect 4863 -288 4879 288
rect 4913 -288 4929 288
rect 4863 -300 4929 -288
rect 4959 288 5025 300
rect 4959 -288 4975 288
rect 5009 -288 5025 288
rect 4959 -300 5025 -288
rect 5055 288 5121 300
rect 5055 -288 5071 288
rect 5105 -288 5121 288
rect 5055 -300 5121 -288
rect 5151 288 5217 300
rect 5151 -288 5167 288
rect 5201 -288 5217 288
rect 5151 -300 5217 -288
rect 5247 288 5313 300
rect 5247 -288 5263 288
rect 5297 -288 5313 288
rect 5247 -300 5313 -288
rect 5343 288 5409 300
rect 5343 -288 5359 288
rect 5393 -288 5409 288
rect 5343 -300 5409 -288
rect 5439 288 5505 300
rect 5439 -288 5455 288
rect 5489 -288 5505 288
rect 5439 -300 5505 -288
rect 5535 288 5601 300
rect 5535 -288 5551 288
rect 5585 -288 5601 288
rect 5535 -300 5601 -288
rect 5631 288 5697 300
rect 5631 -288 5647 288
rect 5681 -288 5697 288
rect 5631 -300 5697 -288
rect 5727 288 5789 300
rect 5727 -288 5743 288
rect 5777 -288 5789 288
rect 5727 -300 5789 -288
<< pdiffc >>
rect -5777 -288 -5743 288
rect -5681 -288 -5647 288
rect -5585 -288 -5551 288
rect -5489 -288 -5455 288
rect -5393 -288 -5359 288
rect -5297 -288 -5263 288
rect -5201 -288 -5167 288
rect -5105 -288 -5071 288
rect -5009 -288 -4975 288
rect -4913 -288 -4879 288
rect -4817 -288 -4783 288
rect -4721 -288 -4687 288
rect -4625 -288 -4591 288
rect -4529 -288 -4495 288
rect -4433 -288 -4399 288
rect -4337 -288 -4303 288
rect -4241 -288 -4207 288
rect -4145 -288 -4111 288
rect -4049 -288 -4015 288
rect -3953 -288 -3919 288
rect -3857 -288 -3823 288
rect -3761 -288 -3727 288
rect -3665 -288 -3631 288
rect -3569 -288 -3535 288
rect -3473 -288 -3439 288
rect -3377 -288 -3343 288
rect -3281 -288 -3247 288
rect -3185 -288 -3151 288
rect -3089 -288 -3055 288
rect -2993 -288 -2959 288
rect -2897 -288 -2863 288
rect -2801 -288 -2767 288
rect -2705 -288 -2671 288
rect -2609 -288 -2575 288
rect -2513 -288 -2479 288
rect -2417 -288 -2383 288
rect -2321 -288 -2287 288
rect -2225 -288 -2191 288
rect -2129 -288 -2095 288
rect -2033 -288 -1999 288
rect -1937 -288 -1903 288
rect -1841 -288 -1807 288
rect -1745 -288 -1711 288
rect -1649 -288 -1615 288
rect -1553 -288 -1519 288
rect -1457 -288 -1423 288
rect -1361 -288 -1327 288
rect -1265 -288 -1231 288
rect -1169 -288 -1135 288
rect -1073 -288 -1039 288
rect -977 -288 -943 288
rect -881 -288 -847 288
rect -785 -288 -751 288
rect -689 -288 -655 288
rect -593 -288 -559 288
rect -497 -288 -463 288
rect -401 -288 -367 288
rect -305 -288 -271 288
rect -209 -288 -175 288
rect -113 -288 -79 288
rect -17 -288 17 288
rect 79 -288 113 288
rect 175 -288 209 288
rect 271 -288 305 288
rect 367 -288 401 288
rect 463 -288 497 288
rect 559 -288 593 288
rect 655 -288 689 288
rect 751 -288 785 288
rect 847 -288 881 288
rect 943 -288 977 288
rect 1039 -288 1073 288
rect 1135 -288 1169 288
rect 1231 -288 1265 288
rect 1327 -288 1361 288
rect 1423 -288 1457 288
rect 1519 -288 1553 288
rect 1615 -288 1649 288
rect 1711 -288 1745 288
rect 1807 -288 1841 288
rect 1903 -288 1937 288
rect 1999 -288 2033 288
rect 2095 -288 2129 288
rect 2191 -288 2225 288
rect 2287 -288 2321 288
rect 2383 -288 2417 288
rect 2479 -288 2513 288
rect 2575 -288 2609 288
rect 2671 -288 2705 288
rect 2767 -288 2801 288
rect 2863 -288 2897 288
rect 2959 -288 2993 288
rect 3055 -288 3089 288
rect 3151 -288 3185 288
rect 3247 -288 3281 288
rect 3343 -288 3377 288
rect 3439 -288 3473 288
rect 3535 -288 3569 288
rect 3631 -288 3665 288
rect 3727 -288 3761 288
rect 3823 -288 3857 288
rect 3919 -288 3953 288
rect 4015 -288 4049 288
rect 4111 -288 4145 288
rect 4207 -288 4241 288
rect 4303 -288 4337 288
rect 4399 -288 4433 288
rect 4495 -288 4529 288
rect 4591 -288 4625 288
rect 4687 -288 4721 288
rect 4783 -288 4817 288
rect 4879 -288 4913 288
rect 4975 -288 5009 288
rect 5071 -288 5105 288
rect 5167 -288 5201 288
rect 5263 -288 5297 288
rect 5359 -288 5393 288
rect 5455 -288 5489 288
rect 5551 -288 5585 288
rect 5647 -288 5681 288
rect 5743 -288 5777 288
<< nsubdiff >>
rect -5891 449 -5795 483
rect 5795 449 5891 483
rect -5891 387 -5857 449
rect 5857 387 5891 449
rect -5891 -449 -5857 -387
rect 5857 -449 5891 -387
rect -5891 -483 -5795 -449
rect 5795 -483 5891 -449
<< nsubdiffcont >>
rect -5795 449 5795 483
rect -5891 -387 -5857 387
rect 5857 -387 5891 387
rect -5795 -483 5795 -449
<< poly >>
rect -5745 381 5745 397
rect -5745 347 -5729 381
rect -5695 347 -5633 381
rect -5599 347 -5537 381
rect -5503 347 -5441 381
rect -5407 347 -5345 381
rect -5311 347 -5249 381
rect -5215 347 -5153 381
rect -5119 347 -5057 381
rect -5023 347 -4961 381
rect -4927 347 -4865 381
rect -4831 347 -4769 381
rect -4735 347 -4673 381
rect -4639 347 -4577 381
rect -4543 347 -4481 381
rect -4447 347 -4385 381
rect -4351 347 -4289 381
rect -4255 347 -4193 381
rect -4159 347 -4097 381
rect -4063 347 -4001 381
rect -3967 347 -3905 381
rect -3871 347 -3809 381
rect -3775 347 -3713 381
rect -3679 347 -3617 381
rect -3583 347 -3521 381
rect -3487 347 -3425 381
rect -3391 347 -3329 381
rect -3295 347 -3233 381
rect -3199 347 -3137 381
rect -3103 347 -3041 381
rect -3007 347 -2945 381
rect -2911 347 -2849 381
rect -2815 347 -2753 381
rect -2719 347 -2657 381
rect -2623 347 -2561 381
rect -2527 347 -2465 381
rect -2431 347 -2369 381
rect -2335 347 -2273 381
rect -2239 347 -2177 381
rect -2143 347 -2081 381
rect -2047 347 -1985 381
rect -1951 347 -1889 381
rect -1855 347 -1793 381
rect -1759 347 -1697 381
rect -1663 347 -1601 381
rect -1567 347 -1505 381
rect -1471 347 -1409 381
rect -1375 347 -1313 381
rect -1279 347 -1217 381
rect -1183 347 -1121 381
rect -1087 347 -1025 381
rect -991 347 -929 381
rect -895 347 -833 381
rect -799 347 -737 381
rect -703 347 -641 381
rect -607 347 -545 381
rect -511 347 -449 381
rect -415 347 -353 381
rect -319 347 -257 381
rect -223 347 -161 381
rect -127 347 -65 381
rect -31 347 31 381
rect 65 347 127 381
rect 161 347 223 381
rect 257 347 319 381
rect 353 347 415 381
rect 449 347 511 381
rect 545 347 607 381
rect 641 347 703 381
rect 737 347 799 381
rect 833 347 895 381
rect 929 347 991 381
rect 1025 347 1087 381
rect 1121 347 1183 381
rect 1217 347 1279 381
rect 1313 347 1375 381
rect 1409 347 1471 381
rect 1505 347 1567 381
rect 1601 347 1663 381
rect 1697 347 1759 381
rect 1793 347 1855 381
rect 1889 347 1951 381
rect 1985 347 2047 381
rect 2081 347 2143 381
rect 2177 347 2239 381
rect 2273 347 2335 381
rect 2369 347 2431 381
rect 2465 347 2527 381
rect 2561 347 2623 381
rect 2657 347 2719 381
rect 2753 347 2815 381
rect 2849 347 2911 381
rect 2945 347 3007 381
rect 3041 347 3103 381
rect 3137 347 3199 381
rect 3233 347 3295 381
rect 3329 347 3391 381
rect 3425 347 3487 381
rect 3521 347 3583 381
rect 3617 347 3679 381
rect 3713 347 3775 381
rect 3809 347 3871 381
rect 3905 347 3967 381
rect 4001 347 4063 381
rect 4097 347 4159 381
rect 4193 347 4255 381
rect 4289 347 4351 381
rect 4385 347 4447 381
rect 4481 347 4543 381
rect 4577 347 4639 381
rect 4673 347 4735 381
rect 4769 347 4831 381
rect 4865 347 4927 381
rect 4961 347 5023 381
rect 5057 347 5119 381
rect 5153 347 5215 381
rect 5249 347 5311 381
rect 5345 347 5407 381
rect 5441 347 5503 381
rect 5537 347 5599 381
rect 5633 347 5695 381
rect 5729 347 5745 381
rect -5745 331 5745 347
rect -5727 300 -5697 331
rect -5631 300 -5601 331
rect -5535 300 -5505 331
rect -5439 300 -5409 331
rect -5343 300 -5313 331
rect -5247 300 -5217 331
rect -5151 300 -5121 331
rect -5055 300 -5025 331
rect -4959 300 -4929 331
rect -4863 300 -4833 331
rect -4767 300 -4737 331
rect -4671 300 -4641 331
rect -4575 300 -4545 331
rect -4479 300 -4449 331
rect -4383 300 -4353 331
rect -4287 300 -4257 331
rect -4191 300 -4161 331
rect -4095 300 -4065 331
rect -3999 300 -3969 331
rect -3903 300 -3873 331
rect -3807 300 -3777 331
rect -3711 300 -3681 331
rect -3615 300 -3585 331
rect -3519 300 -3489 331
rect -3423 300 -3393 331
rect -3327 300 -3297 331
rect -3231 300 -3201 331
rect -3135 300 -3105 331
rect -3039 300 -3009 331
rect -2943 300 -2913 331
rect -2847 300 -2817 331
rect -2751 300 -2721 331
rect -2655 300 -2625 331
rect -2559 300 -2529 331
rect -2463 300 -2433 331
rect -2367 300 -2337 331
rect -2271 300 -2241 331
rect -2175 300 -2145 331
rect -2079 300 -2049 331
rect -1983 300 -1953 331
rect -1887 300 -1857 331
rect -1791 300 -1761 331
rect -1695 300 -1665 331
rect -1599 300 -1569 331
rect -1503 300 -1473 331
rect -1407 300 -1377 331
rect -1311 300 -1281 331
rect -1215 300 -1185 331
rect -1119 300 -1089 331
rect -1023 300 -993 331
rect -927 300 -897 331
rect -831 300 -801 331
rect -735 300 -705 331
rect -639 300 -609 331
rect -543 300 -513 331
rect -447 300 -417 331
rect -351 300 -321 331
rect -255 300 -225 331
rect -159 300 -129 331
rect -63 300 -33 331
rect 33 300 63 331
rect 129 300 159 331
rect 225 300 255 331
rect 321 300 351 331
rect 417 300 447 331
rect 513 300 543 331
rect 609 300 639 331
rect 705 300 735 331
rect 801 300 831 331
rect 897 300 927 331
rect 993 300 1023 331
rect 1089 300 1119 331
rect 1185 300 1215 331
rect 1281 300 1311 331
rect 1377 300 1407 331
rect 1473 300 1503 331
rect 1569 300 1599 331
rect 1665 300 1695 331
rect 1761 300 1791 331
rect 1857 300 1887 331
rect 1953 300 1983 331
rect 2049 300 2079 331
rect 2145 300 2175 331
rect 2241 300 2271 331
rect 2337 300 2367 331
rect 2433 300 2463 331
rect 2529 300 2559 331
rect 2625 300 2655 331
rect 2721 300 2751 331
rect 2817 300 2847 331
rect 2913 300 2943 331
rect 3009 300 3039 331
rect 3105 300 3135 331
rect 3201 300 3231 331
rect 3297 300 3327 331
rect 3393 300 3423 331
rect 3489 300 3519 331
rect 3585 300 3615 331
rect 3681 300 3711 331
rect 3777 300 3807 331
rect 3873 300 3903 331
rect 3969 300 3999 331
rect 4065 300 4095 331
rect 4161 300 4191 331
rect 4257 300 4287 331
rect 4353 300 4383 331
rect 4449 300 4479 331
rect 4545 300 4575 331
rect 4641 300 4671 331
rect 4737 300 4767 331
rect 4833 300 4863 331
rect 4929 300 4959 331
rect 5025 300 5055 331
rect 5121 300 5151 331
rect 5217 300 5247 331
rect 5313 300 5343 331
rect 5409 300 5439 331
rect 5505 300 5535 331
rect 5601 300 5631 331
rect 5697 300 5727 331
rect -5727 -331 -5697 -300
rect -5631 -331 -5601 -300
rect -5535 -331 -5505 -300
rect -5439 -331 -5409 -300
rect -5343 -331 -5313 -300
rect -5247 -331 -5217 -300
rect -5151 -331 -5121 -300
rect -5055 -331 -5025 -300
rect -4959 -331 -4929 -300
rect -4863 -331 -4833 -300
rect -4767 -331 -4737 -300
rect -4671 -331 -4641 -300
rect -4575 -331 -4545 -300
rect -4479 -331 -4449 -300
rect -4383 -331 -4353 -300
rect -4287 -331 -4257 -300
rect -4191 -331 -4161 -300
rect -4095 -331 -4065 -300
rect -3999 -331 -3969 -300
rect -3903 -331 -3873 -300
rect -3807 -331 -3777 -300
rect -3711 -331 -3681 -300
rect -3615 -331 -3585 -300
rect -3519 -331 -3489 -300
rect -3423 -331 -3393 -300
rect -3327 -331 -3297 -300
rect -3231 -331 -3201 -300
rect -3135 -331 -3105 -300
rect -3039 -331 -3009 -300
rect -2943 -331 -2913 -300
rect -2847 -331 -2817 -300
rect -2751 -331 -2721 -300
rect -2655 -331 -2625 -300
rect -2559 -331 -2529 -300
rect -2463 -331 -2433 -300
rect -2367 -331 -2337 -300
rect -2271 -331 -2241 -300
rect -2175 -331 -2145 -300
rect -2079 -331 -2049 -300
rect -1983 -331 -1953 -300
rect -1887 -331 -1857 -300
rect -1791 -331 -1761 -300
rect -1695 -331 -1665 -300
rect -1599 -331 -1569 -300
rect -1503 -331 -1473 -300
rect -1407 -331 -1377 -300
rect -1311 -331 -1281 -300
rect -1215 -331 -1185 -300
rect -1119 -331 -1089 -300
rect -1023 -331 -993 -300
rect -927 -331 -897 -300
rect -831 -331 -801 -300
rect -735 -331 -705 -300
rect -639 -331 -609 -300
rect -543 -331 -513 -300
rect -447 -331 -417 -300
rect -351 -331 -321 -300
rect -255 -331 -225 -300
rect -159 -331 -129 -300
rect -63 -331 -33 -300
rect 33 -331 63 -300
rect 129 -331 159 -300
rect 225 -331 255 -300
rect 321 -331 351 -300
rect 417 -331 447 -300
rect 513 -331 543 -300
rect 609 -331 639 -300
rect 705 -331 735 -300
rect 801 -331 831 -300
rect 897 -331 927 -300
rect 993 -331 1023 -300
rect 1089 -331 1119 -300
rect 1185 -331 1215 -300
rect 1281 -331 1311 -300
rect 1377 -331 1407 -300
rect 1473 -331 1503 -300
rect 1569 -331 1599 -300
rect 1665 -331 1695 -300
rect 1761 -331 1791 -300
rect 1857 -331 1887 -300
rect 1953 -331 1983 -300
rect 2049 -331 2079 -300
rect 2145 -331 2175 -300
rect 2241 -331 2271 -300
rect 2337 -331 2367 -300
rect 2433 -331 2463 -300
rect 2529 -331 2559 -300
rect 2625 -331 2655 -300
rect 2721 -331 2751 -300
rect 2817 -331 2847 -300
rect 2913 -331 2943 -300
rect 3009 -331 3039 -300
rect 3105 -331 3135 -300
rect 3201 -331 3231 -300
rect 3297 -331 3327 -300
rect 3393 -331 3423 -300
rect 3489 -331 3519 -300
rect 3585 -331 3615 -300
rect 3681 -331 3711 -300
rect 3777 -331 3807 -300
rect 3873 -331 3903 -300
rect 3969 -331 3999 -300
rect 4065 -331 4095 -300
rect 4161 -331 4191 -300
rect 4257 -331 4287 -300
rect 4353 -331 4383 -300
rect 4449 -331 4479 -300
rect 4545 -331 4575 -300
rect 4641 -331 4671 -300
rect 4737 -331 4767 -300
rect 4833 -331 4863 -300
rect 4929 -331 4959 -300
rect 5025 -331 5055 -300
rect 5121 -331 5151 -300
rect 5217 -331 5247 -300
rect 5313 -331 5343 -300
rect 5409 -331 5439 -300
rect 5505 -331 5535 -300
rect 5601 -331 5631 -300
rect 5697 -331 5727 -300
rect -5745 -347 5745 -331
rect -5745 -381 -5729 -347
rect -5695 -381 -5633 -347
rect -5599 -381 -5537 -347
rect -5503 -381 -5441 -347
rect -5407 -381 -5345 -347
rect -5311 -381 -5249 -347
rect -5215 -381 -5153 -347
rect -5119 -381 -5057 -347
rect -5023 -381 -4961 -347
rect -4927 -381 -4865 -347
rect -4831 -381 -4769 -347
rect -4735 -381 -4673 -347
rect -4639 -381 -4577 -347
rect -4543 -381 -4481 -347
rect -4447 -381 -4385 -347
rect -4351 -381 -4289 -347
rect -4255 -381 -4193 -347
rect -4159 -381 -4097 -347
rect -4063 -381 -4001 -347
rect -3967 -381 -3905 -347
rect -3871 -381 -3809 -347
rect -3775 -381 -3713 -347
rect -3679 -381 -3617 -347
rect -3583 -381 -3521 -347
rect -3487 -381 -3425 -347
rect -3391 -381 -3329 -347
rect -3295 -381 -3233 -347
rect -3199 -381 -3137 -347
rect -3103 -381 -3041 -347
rect -3007 -381 -2945 -347
rect -2911 -381 -2849 -347
rect -2815 -381 -2753 -347
rect -2719 -381 -2657 -347
rect -2623 -381 -2561 -347
rect -2527 -381 -2465 -347
rect -2431 -381 -2369 -347
rect -2335 -381 -2273 -347
rect -2239 -381 -2177 -347
rect -2143 -381 -2081 -347
rect -2047 -381 -1985 -347
rect -1951 -381 -1889 -347
rect -1855 -381 -1793 -347
rect -1759 -381 -1697 -347
rect -1663 -381 -1601 -347
rect -1567 -381 -1505 -347
rect -1471 -381 -1409 -347
rect -1375 -381 -1313 -347
rect -1279 -381 -1217 -347
rect -1183 -381 -1121 -347
rect -1087 -381 -1025 -347
rect -991 -381 -929 -347
rect -895 -381 -833 -347
rect -799 -381 -737 -347
rect -703 -381 -641 -347
rect -607 -381 -545 -347
rect -511 -381 -449 -347
rect -415 -381 -353 -347
rect -319 -381 -257 -347
rect -223 -381 -161 -347
rect -127 -381 -65 -347
rect -31 -381 31 -347
rect 65 -381 127 -347
rect 161 -381 223 -347
rect 257 -381 319 -347
rect 353 -381 415 -347
rect 449 -381 511 -347
rect 545 -381 607 -347
rect 641 -381 703 -347
rect 737 -381 799 -347
rect 833 -381 895 -347
rect 929 -381 991 -347
rect 1025 -381 1087 -347
rect 1121 -381 1183 -347
rect 1217 -381 1279 -347
rect 1313 -381 1375 -347
rect 1409 -381 1471 -347
rect 1505 -381 1567 -347
rect 1601 -381 1663 -347
rect 1697 -381 1759 -347
rect 1793 -381 1855 -347
rect 1889 -381 1951 -347
rect 1985 -381 2047 -347
rect 2081 -381 2143 -347
rect 2177 -381 2239 -347
rect 2273 -381 2335 -347
rect 2369 -381 2431 -347
rect 2465 -381 2527 -347
rect 2561 -381 2623 -347
rect 2657 -381 2719 -347
rect 2753 -381 2815 -347
rect 2849 -381 2911 -347
rect 2945 -381 3007 -347
rect 3041 -381 3103 -347
rect 3137 -381 3199 -347
rect 3233 -381 3295 -347
rect 3329 -381 3391 -347
rect 3425 -381 3487 -347
rect 3521 -381 3583 -347
rect 3617 -381 3679 -347
rect 3713 -381 3775 -347
rect 3809 -381 3871 -347
rect 3905 -381 3967 -347
rect 4001 -381 4063 -347
rect 4097 -381 4159 -347
rect 4193 -381 4255 -347
rect 4289 -381 4351 -347
rect 4385 -381 4447 -347
rect 4481 -381 4543 -347
rect 4577 -381 4639 -347
rect 4673 -381 4735 -347
rect 4769 -381 4831 -347
rect 4865 -381 4927 -347
rect 4961 -381 5023 -347
rect 5057 -381 5119 -347
rect 5153 -381 5215 -347
rect 5249 -381 5311 -347
rect 5345 -381 5407 -347
rect 5441 -381 5503 -347
rect 5537 -381 5599 -347
rect 5633 -381 5695 -347
rect 5729 -381 5745 -347
rect -5745 -397 5745 -381
<< polycont >>
rect -5729 347 -5695 381
rect -5633 347 -5599 381
rect -5537 347 -5503 381
rect -5441 347 -5407 381
rect -5345 347 -5311 381
rect -5249 347 -5215 381
rect -5153 347 -5119 381
rect -5057 347 -5023 381
rect -4961 347 -4927 381
rect -4865 347 -4831 381
rect -4769 347 -4735 381
rect -4673 347 -4639 381
rect -4577 347 -4543 381
rect -4481 347 -4447 381
rect -4385 347 -4351 381
rect -4289 347 -4255 381
rect -4193 347 -4159 381
rect -4097 347 -4063 381
rect -4001 347 -3967 381
rect -3905 347 -3871 381
rect -3809 347 -3775 381
rect -3713 347 -3679 381
rect -3617 347 -3583 381
rect -3521 347 -3487 381
rect -3425 347 -3391 381
rect -3329 347 -3295 381
rect -3233 347 -3199 381
rect -3137 347 -3103 381
rect -3041 347 -3007 381
rect -2945 347 -2911 381
rect -2849 347 -2815 381
rect -2753 347 -2719 381
rect -2657 347 -2623 381
rect -2561 347 -2527 381
rect -2465 347 -2431 381
rect -2369 347 -2335 381
rect -2273 347 -2239 381
rect -2177 347 -2143 381
rect -2081 347 -2047 381
rect -1985 347 -1951 381
rect -1889 347 -1855 381
rect -1793 347 -1759 381
rect -1697 347 -1663 381
rect -1601 347 -1567 381
rect -1505 347 -1471 381
rect -1409 347 -1375 381
rect -1313 347 -1279 381
rect -1217 347 -1183 381
rect -1121 347 -1087 381
rect -1025 347 -991 381
rect -929 347 -895 381
rect -833 347 -799 381
rect -737 347 -703 381
rect -641 347 -607 381
rect -545 347 -511 381
rect -449 347 -415 381
rect -353 347 -319 381
rect -257 347 -223 381
rect -161 347 -127 381
rect -65 347 -31 381
rect 31 347 65 381
rect 127 347 161 381
rect 223 347 257 381
rect 319 347 353 381
rect 415 347 449 381
rect 511 347 545 381
rect 607 347 641 381
rect 703 347 737 381
rect 799 347 833 381
rect 895 347 929 381
rect 991 347 1025 381
rect 1087 347 1121 381
rect 1183 347 1217 381
rect 1279 347 1313 381
rect 1375 347 1409 381
rect 1471 347 1505 381
rect 1567 347 1601 381
rect 1663 347 1697 381
rect 1759 347 1793 381
rect 1855 347 1889 381
rect 1951 347 1985 381
rect 2047 347 2081 381
rect 2143 347 2177 381
rect 2239 347 2273 381
rect 2335 347 2369 381
rect 2431 347 2465 381
rect 2527 347 2561 381
rect 2623 347 2657 381
rect 2719 347 2753 381
rect 2815 347 2849 381
rect 2911 347 2945 381
rect 3007 347 3041 381
rect 3103 347 3137 381
rect 3199 347 3233 381
rect 3295 347 3329 381
rect 3391 347 3425 381
rect 3487 347 3521 381
rect 3583 347 3617 381
rect 3679 347 3713 381
rect 3775 347 3809 381
rect 3871 347 3905 381
rect 3967 347 4001 381
rect 4063 347 4097 381
rect 4159 347 4193 381
rect 4255 347 4289 381
rect 4351 347 4385 381
rect 4447 347 4481 381
rect 4543 347 4577 381
rect 4639 347 4673 381
rect 4735 347 4769 381
rect 4831 347 4865 381
rect 4927 347 4961 381
rect 5023 347 5057 381
rect 5119 347 5153 381
rect 5215 347 5249 381
rect 5311 347 5345 381
rect 5407 347 5441 381
rect 5503 347 5537 381
rect 5599 347 5633 381
rect 5695 347 5729 381
rect -5729 -381 -5695 -347
rect -5633 -381 -5599 -347
rect -5537 -381 -5503 -347
rect -5441 -381 -5407 -347
rect -5345 -381 -5311 -347
rect -5249 -381 -5215 -347
rect -5153 -381 -5119 -347
rect -5057 -381 -5023 -347
rect -4961 -381 -4927 -347
rect -4865 -381 -4831 -347
rect -4769 -381 -4735 -347
rect -4673 -381 -4639 -347
rect -4577 -381 -4543 -347
rect -4481 -381 -4447 -347
rect -4385 -381 -4351 -347
rect -4289 -381 -4255 -347
rect -4193 -381 -4159 -347
rect -4097 -381 -4063 -347
rect -4001 -381 -3967 -347
rect -3905 -381 -3871 -347
rect -3809 -381 -3775 -347
rect -3713 -381 -3679 -347
rect -3617 -381 -3583 -347
rect -3521 -381 -3487 -347
rect -3425 -381 -3391 -347
rect -3329 -381 -3295 -347
rect -3233 -381 -3199 -347
rect -3137 -381 -3103 -347
rect -3041 -381 -3007 -347
rect -2945 -381 -2911 -347
rect -2849 -381 -2815 -347
rect -2753 -381 -2719 -347
rect -2657 -381 -2623 -347
rect -2561 -381 -2527 -347
rect -2465 -381 -2431 -347
rect -2369 -381 -2335 -347
rect -2273 -381 -2239 -347
rect -2177 -381 -2143 -347
rect -2081 -381 -2047 -347
rect -1985 -381 -1951 -347
rect -1889 -381 -1855 -347
rect -1793 -381 -1759 -347
rect -1697 -381 -1663 -347
rect -1601 -381 -1567 -347
rect -1505 -381 -1471 -347
rect -1409 -381 -1375 -347
rect -1313 -381 -1279 -347
rect -1217 -381 -1183 -347
rect -1121 -381 -1087 -347
rect -1025 -381 -991 -347
rect -929 -381 -895 -347
rect -833 -381 -799 -347
rect -737 -381 -703 -347
rect -641 -381 -607 -347
rect -545 -381 -511 -347
rect -449 -381 -415 -347
rect -353 -381 -319 -347
rect -257 -381 -223 -347
rect -161 -381 -127 -347
rect -65 -381 -31 -347
rect 31 -381 65 -347
rect 127 -381 161 -347
rect 223 -381 257 -347
rect 319 -381 353 -347
rect 415 -381 449 -347
rect 511 -381 545 -347
rect 607 -381 641 -347
rect 703 -381 737 -347
rect 799 -381 833 -347
rect 895 -381 929 -347
rect 991 -381 1025 -347
rect 1087 -381 1121 -347
rect 1183 -381 1217 -347
rect 1279 -381 1313 -347
rect 1375 -381 1409 -347
rect 1471 -381 1505 -347
rect 1567 -381 1601 -347
rect 1663 -381 1697 -347
rect 1759 -381 1793 -347
rect 1855 -381 1889 -347
rect 1951 -381 1985 -347
rect 2047 -381 2081 -347
rect 2143 -381 2177 -347
rect 2239 -381 2273 -347
rect 2335 -381 2369 -347
rect 2431 -381 2465 -347
rect 2527 -381 2561 -347
rect 2623 -381 2657 -347
rect 2719 -381 2753 -347
rect 2815 -381 2849 -347
rect 2911 -381 2945 -347
rect 3007 -381 3041 -347
rect 3103 -381 3137 -347
rect 3199 -381 3233 -347
rect 3295 -381 3329 -347
rect 3391 -381 3425 -347
rect 3487 -381 3521 -347
rect 3583 -381 3617 -347
rect 3679 -381 3713 -347
rect 3775 -381 3809 -347
rect 3871 -381 3905 -347
rect 3967 -381 4001 -347
rect 4063 -381 4097 -347
rect 4159 -381 4193 -347
rect 4255 -381 4289 -347
rect 4351 -381 4385 -347
rect 4447 -381 4481 -347
rect 4543 -381 4577 -347
rect 4639 -381 4673 -347
rect 4735 -381 4769 -347
rect 4831 -381 4865 -347
rect 4927 -381 4961 -347
rect 5023 -381 5057 -347
rect 5119 -381 5153 -347
rect 5215 -381 5249 -347
rect 5311 -381 5345 -347
rect 5407 -381 5441 -347
rect 5503 -381 5537 -347
rect 5599 -381 5633 -347
rect 5695 -381 5729 -347
<< locali >>
rect -5891 449 -5885 483
rect 5795 449 5891 483
rect -5891 387 -5857 449
rect 5857 387 5891 449
rect -5745 347 -5729 381
rect -5695 347 -5633 381
rect -5599 347 -5537 381
rect -5503 347 -5441 381
rect -5407 347 -5345 381
rect -5311 347 -5249 381
rect -5215 347 -5153 381
rect -5119 347 -5057 381
rect -5023 347 -4961 381
rect -4927 347 -4865 381
rect -4831 347 -4769 381
rect -4735 347 -4673 381
rect -4639 347 -4577 381
rect -4543 347 -4481 381
rect -4447 347 -4385 381
rect -4351 347 -4289 381
rect -4255 347 -4193 381
rect -4159 347 -4097 381
rect -4063 347 -4001 381
rect -3967 347 -3905 381
rect -3871 347 -3809 381
rect -3775 347 -3713 381
rect -3679 347 -3617 381
rect -3583 347 -3521 381
rect -3487 347 -3425 381
rect -3391 347 -3329 381
rect -3295 347 -3233 381
rect -3199 347 -3137 381
rect -3103 347 -3041 381
rect -3007 347 -2945 381
rect -2911 347 -2849 381
rect -2815 347 -2753 381
rect -2719 347 -2657 381
rect -2623 347 -2561 381
rect -2527 347 -2465 381
rect -2431 347 -2369 381
rect -2335 347 -2273 381
rect -2239 347 -2177 381
rect -2143 347 -2081 381
rect -2047 347 -1985 381
rect -1951 347 -1889 381
rect -1855 347 -1793 381
rect -1759 347 -1697 381
rect -1663 347 -1601 381
rect -1567 347 -1505 381
rect -1471 347 -1409 381
rect -1375 347 -1313 381
rect -1279 347 -1217 381
rect -1183 347 -1121 381
rect -1087 347 -1025 381
rect -991 347 -929 381
rect -895 347 -833 381
rect -799 347 -737 381
rect -703 347 -641 381
rect -607 347 -545 381
rect -511 347 -449 381
rect -415 347 -353 381
rect -319 347 -257 381
rect -223 347 -161 381
rect -127 347 -65 381
rect -31 347 31 381
rect 65 347 127 381
rect 161 347 223 381
rect 257 347 319 381
rect 353 347 415 381
rect 449 347 511 381
rect 545 347 607 381
rect 641 347 703 381
rect 737 347 799 381
rect 833 347 895 381
rect 929 347 991 381
rect 1025 347 1087 381
rect 1121 347 1183 381
rect 1217 347 1279 381
rect 1313 347 1375 381
rect 1409 347 1471 381
rect 1505 347 1567 381
rect 1601 347 1663 381
rect 1697 347 1759 381
rect 1793 347 1855 381
rect 1889 347 1951 381
rect 1985 347 2047 381
rect 2081 347 2143 381
rect 2177 347 2239 381
rect 2273 347 2335 381
rect 2369 347 2431 381
rect 2465 347 2527 381
rect 2561 347 2623 381
rect 2657 347 2719 381
rect 2753 347 2815 381
rect 2849 347 2911 381
rect 2945 347 3007 381
rect 3041 347 3103 381
rect 3137 347 3199 381
rect 3233 347 3295 381
rect 3329 347 3391 381
rect 3425 347 3487 381
rect 3521 347 3583 381
rect 3617 347 3679 381
rect 3713 347 3775 381
rect 3809 347 3871 381
rect 3905 347 3967 381
rect 4001 347 4063 381
rect 4097 347 4159 381
rect 4193 347 4255 381
rect 4289 347 4351 381
rect 4385 347 4447 381
rect 4481 347 4543 381
rect 4577 347 4639 381
rect 4673 347 4735 381
rect 4769 347 4831 381
rect 4865 347 4927 381
rect 4961 347 5023 381
rect 5057 347 5119 381
rect 5153 347 5215 381
rect 5249 347 5311 381
rect 5345 347 5407 381
rect 5441 347 5503 381
rect 5537 347 5599 381
rect 5633 347 5695 381
rect 5729 347 5745 381
rect -5777 288 -5743 304
rect -5777 -304 -5743 -288
rect -5681 288 -5647 304
rect -5681 -304 -5647 -288
rect -5585 288 -5551 304
rect -5585 -304 -5551 -288
rect -5489 288 -5455 304
rect -5489 -304 -5455 -288
rect -5393 288 -5359 304
rect -5393 -304 -5359 -288
rect -5297 288 -5263 304
rect -5297 -304 -5263 -288
rect -5201 288 -5167 304
rect -5201 -304 -5167 -288
rect -5105 288 -5071 304
rect -5105 -304 -5071 -288
rect -5009 288 -4975 304
rect -5009 -304 -4975 -288
rect -4913 288 -4879 304
rect -4913 -304 -4879 -288
rect -4817 288 -4783 304
rect -4817 -304 -4783 -288
rect -4721 288 -4687 304
rect -4721 -304 -4687 -288
rect -4625 288 -4591 304
rect -4625 -304 -4591 -288
rect -4529 288 -4495 304
rect -4529 -304 -4495 -288
rect -4433 288 -4399 304
rect -4433 -304 -4399 -288
rect -4337 288 -4303 304
rect -4337 -304 -4303 -288
rect -4241 288 -4207 304
rect -4241 -304 -4207 -288
rect -4145 288 -4111 304
rect -4145 -304 -4111 -288
rect -4049 288 -4015 304
rect -4049 -304 -4015 -288
rect -3953 288 -3919 304
rect -3953 -304 -3919 -288
rect -3857 288 -3823 304
rect -3857 -304 -3823 -288
rect -3761 288 -3727 304
rect -3761 -304 -3727 -288
rect -3665 288 -3631 304
rect -3665 -304 -3631 -288
rect -3569 288 -3535 304
rect -3569 -304 -3535 -288
rect -3473 288 -3439 304
rect -3473 -304 -3439 -288
rect -3377 288 -3343 304
rect -3377 -304 -3343 -288
rect -3281 288 -3247 304
rect -3281 -304 -3247 -288
rect -3185 288 -3151 304
rect -3185 -304 -3151 -288
rect -3089 288 -3055 304
rect -3089 -304 -3055 -288
rect -2993 288 -2959 304
rect -2993 -304 -2959 -288
rect -2897 288 -2863 304
rect -2897 -304 -2863 -288
rect -2801 288 -2767 304
rect -2801 -304 -2767 -288
rect -2705 288 -2671 304
rect -2705 -304 -2671 -288
rect -2609 288 -2575 304
rect -2609 -304 -2575 -288
rect -2513 288 -2479 304
rect -2513 -304 -2479 -288
rect -2417 288 -2383 304
rect -2417 -304 -2383 -288
rect -2321 288 -2287 304
rect -2321 -304 -2287 -288
rect -2225 288 -2191 304
rect -2225 -304 -2191 -288
rect -2129 288 -2095 304
rect -2129 -304 -2095 -288
rect -2033 288 -1999 304
rect -2033 -304 -1999 -288
rect -1937 288 -1903 304
rect -1937 -304 -1903 -288
rect -1841 288 -1807 304
rect -1841 -304 -1807 -288
rect -1745 288 -1711 304
rect -1745 -304 -1711 -288
rect -1649 288 -1615 304
rect -1649 -304 -1615 -288
rect -1553 288 -1519 304
rect -1553 -304 -1519 -288
rect -1457 288 -1423 304
rect -1457 -304 -1423 -288
rect -1361 288 -1327 304
rect -1361 -304 -1327 -288
rect -1265 288 -1231 304
rect -1265 -304 -1231 -288
rect -1169 288 -1135 304
rect -1169 -304 -1135 -288
rect -1073 288 -1039 304
rect -1073 -304 -1039 -288
rect -977 288 -943 304
rect -977 -304 -943 -288
rect -881 288 -847 304
rect -881 -304 -847 -288
rect -785 288 -751 304
rect -785 -304 -751 -288
rect -689 288 -655 304
rect -689 -304 -655 -288
rect -593 288 -559 304
rect -593 -304 -559 -288
rect -497 288 -463 304
rect -497 -304 -463 -288
rect -401 288 -367 304
rect -401 -304 -367 -288
rect -305 288 -271 304
rect -305 -304 -271 -288
rect -209 288 -175 304
rect -209 -304 -175 -288
rect -113 288 -79 304
rect -113 -304 -79 -288
rect -17 288 17 304
rect -17 -304 17 -288
rect 79 288 113 304
rect 79 -304 113 -288
rect 175 288 209 304
rect 175 -304 209 -288
rect 271 288 305 304
rect 271 -304 305 -288
rect 367 288 401 304
rect 367 -304 401 -288
rect 463 288 497 304
rect 463 -304 497 -288
rect 559 288 593 304
rect 559 -304 593 -288
rect 655 288 689 304
rect 655 -304 689 -288
rect 751 288 785 304
rect 751 -304 785 -288
rect 847 288 881 304
rect 847 -304 881 -288
rect 943 288 977 304
rect 943 -304 977 -288
rect 1039 288 1073 304
rect 1039 -304 1073 -288
rect 1135 288 1169 304
rect 1135 -304 1169 -288
rect 1231 288 1265 304
rect 1231 -304 1265 -288
rect 1327 288 1361 304
rect 1327 -304 1361 -288
rect 1423 288 1457 304
rect 1423 -304 1457 -288
rect 1519 288 1553 304
rect 1519 -304 1553 -288
rect 1615 288 1649 304
rect 1615 -304 1649 -288
rect 1711 288 1745 304
rect 1711 -304 1745 -288
rect 1807 288 1841 304
rect 1807 -304 1841 -288
rect 1903 288 1937 304
rect 1903 -304 1937 -288
rect 1999 288 2033 304
rect 1999 -304 2033 -288
rect 2095 288 2129 304
rect 2095 -304 2129 -288
rect 2191 288 2225 304
rect 2191 -304 2225 -288
rect 2287 288 2321 304
rect 2287 -304 2321 -288
rect 2383 288 2417 304
rect 2383 -304 2417 -288
rect 2479 288 2513 304
rect 2479 -304 2513 -288
rect 2575 288 2609 304
rect 2575 -304 2609 -288
rect 2671 288 2705 304
rect 2671 -304 2705 -288
rect 2767 288 2801 304
rect 2767 -304 2801 -288
rect 2863 288 2897 304
rect 2863 -304 2897 -288
rect 2959 288 2993 304
rect 2959 -304 2993 -288
rect 3055 288 3089 304
rect 3055 -304 3089 -288
rect 3151 288 3185 304
rect 3151 -304 3185 -288
rect 3247 288 3281 304
rect 3247 -304 3281 -288
rect 3343 288 3377 304
rect 3343 -304 3377 -288
rect 3439 288 3473 304
rect 3439 -304 3473 -288
rect 3535 288 3569 304
rect 3535 -304 3569 -288
rect 3631 288 3665 304
rect 3631 -304 3665 -288
rect 3727 288 3761 304
rect 3727 -304 3761 -288
rect 3823 288 3857 304
rect 3823 -304 3857 -288
rect 3919 288 3953 304
rect 3919 -304 3953 -288
rect 4015 288 4049 304
rect 4015 -304 4049 -288
rect 4111 288 4145 304
rect 4111 -304 4145 -288
rect 4207 288 4241 304
rect 4207 -304 4241 -288
rect 4303 288 4337 304
rect 4303 -304 4337 -288
rect 4399 288 4433 304
rect 4399 -304 4433 -288
rect 4495 288 4529 304
rect 4495 -304 4529 -288
rect 4591 288 4625 304
rect 4591 -304 4625 -288
rect 4687 288 4721 304
rect 4687 -304 4721 -288
rect 4783 288 4817 304
rect 4783 -304 4817 -288
rect 4879 288 4913 304
rect 4879 -304 4913 -288
rect 4975 288 5009 304
rect 4975 -304 5009 -288
rect 5071 288 5105 304
rect 5071 -304 5105 -288
rect 5167 288 5201 304
rect 5167 -304 5201 -288
rect 5263 288 5297 304
rect 5263 -304 5297 -288
rect 5359 288 5393 304
rect 5359 -304 5393 -288
rect 5455 288 5489 304
rect 5455 -304 5489 -288
rect 5551 288 5585 304
rect 5551 -304 5585 -288
rect 5647 288 5681 304
rect 5647 -304 5681 -288
rect 5743 288 5777 304
rect 5743 -304 5777 -288
rect -5745 -381 -5729 -347
rect -5695 -381 -5633 -347
rect -5599 -381 -5537 -347
rect -5503 -381 -5441 -347
rect -5407 -381 -5345 -347
rect -5311 -381 -5249 -347
rect -5215 -381 -5153 -347
rect -5119 -381 -5057 -347
rect -5023 -381 -4961 -347
rect -4927 -381 -4865 -347
rect -4831 -381 -4769 -347
rect -4735 -381 -4673 -347
rect -4639 -381 -4577 -347
rect -4543 -381 -4481 -347
rect -4447 -381 -4385 -347
rect -4351 -381 -4289 -347
rect -4255 -381 -4193 -347
rect -4159 -381 -4097 -347
rect -4063 -381 -4001 -347
rect -3967 -381 -3905 -347
rect -3871 -381 -3809 -347
rect -3775 -381 -3713 -347
rect -3679 -381 -3617 -347
rect -3583 -381 -3521 -347
rect -3487 -381 -3425 -347
rect -3391 -381 -3329 -347
rect -3295 -381 -3233 -347
rect -3199 -381 -3137 -347
rect -3103 -381 -3041 -347
rect -3007 -381 -2945 -347
rect -2911 -381 -2849 -347
rect -2815 -381 -2753 -347
rect -2719 -381 -2657 -347
rect -2623 -381 -2561 -347
rect -2527 -381 -2465 -347
rect -2431 -381 -2369 -347
rect -2335 -381 -2273 -347
rect -2239 -381 -2177 -347
rect -2143 -381 -2081 -347
rect -2047 -381 -1985 -347
rect -1951 -381 -1889 -347
rect -1855 -381 -1793 -347
rect -1759 -381 -1697 -347
rect -1663 -381 -1601 -347
rect -1567 -381 -1505 -347
rect -1471 -381 -1409 -347
rect -1375 -381 -1313 -347
rect -1279 -381 -1217 -347
rect -1183 -381 -1121 -347
rect -1087 -381 -1025 -347
rect -991 -381 -929 -347
rect -895 -381 -833 -347
rect -799 -381 -737 -347
rect -703 -381 -641 -347
rect -607 -381 -545 -347
rect -511 -381 -449 -347
rect -415 -381 -353 -347
rect -319 -381 -257 -347
rect -223 -381 -161 -347
rect -127 -381 -65 -347
rect -31 -381 31 -347
rect 65 -381 127 -347
rect 161 -381 223 -347
rect 257 -381 319 -347
rect 353 -381 415 -347
rect 449 -381 511 -347
rect 545 -381 607 -347
rect 641 -381 703 -347
rect 737 -381 799 -347
rect 833 -381 895 -347
rect 929 -381 991 -347
rect 1025 -381 1087 -347
rect 1121 -381 1183 -347
rect 1217 -381 1279 -347
rect 1313 -381 1375 -347
rect 1409 -381 1471 -347
rect 1505 -381 1567 -347
rect 1601 -381 1663 -347
rect 1697 -381 1759 -347
rect 1793 -381 1855 -347
rect 1889 -381 1951 -347
rect 1985 -381 2047 -347
rect 2081 -381 2143 -347
rect 2177 -381 2239 -347
rect 2273 -381 2335 -347
rect 2369 -381 2431 -347
rect 2465 -381 2527 -347
rect 2561 -381 2623 -347
rect 2657 -381 2719 -347
rect 2753 -381 2815 -347
rect 2849 -381 2911 -347
rect 2945 -381 3007 -347
rect 3041 -381 3103 -347
rect 3137 -381 3199 -347
rect 3233 -381 3295 -347
rect 3329 -381 3391 -347
rect 3425 -381 3487 -347
rect 3521 -381 3583 -347
rect 3617 -381 3679 -347
rect 3713 -381 3775 -347
rect 3809 -381 3871 -347
rect 3905 -381 3967 -347
rect 4001 -381 4063 -347
rect 4097 -381 4159 -347
rect 4193 -381 4255 -347
rect 4289 -381 4351 -347
rect 4385 -381 4447 -347
rect 4481 -381 4543 -347
rect 4577 -381 4639 -347
rect 4673 -381 4735 -347
rect 4769 -381 4831 -347
rect 4865 -381 4927 -347
rect 4961 -381 5023 -347
rect 5057 -381 5119 -347
rect 5153 -381 5215 -347
rect 5249 -381 5311 -347
rect 5345 -381 5407 -347
rect 5441 -381 5503 -347
rect 5537 -381 5599 -347
rect 5633 -381 5695 -347
rect 5729 -381 5745 -347
rect -5891 -449 -5857 -387
rect 5857 -449 5891 -387
rect -5891 -483 -5885 -449
rect 5795 -483 5891 -449
<< viali >>
rect -5885 449 -5795 483
rect -5795 449 5795 483
rect -5729 347 -5695 381
rect -5633 347 -5599 381
rect -5537 347 -5503 381
rect -5441 347 -5407 381
rect -5345 347 -5311 381
rect -5249 347 -5215 381
rect -5153 347 -5119 381
rect -5057 347 -5023 381
rect -4961 347 -4927 381
rect -4865 347 -4831 381
rect -4769 347 -4735 381
rect -4673 347 -4639 381
rect -4577 347 -4543 381
rect -4481 347 -4447 381
rect -4385 347 -4351 381
rect -4289 347 -4255 381
rect -4193 347 -4159 381
rect -4097 347 -4063 381
rect -4001 347 -3967 381
rect -3905 347 -3871 381
rect -3809 347 -3775 381
rect -3713 347 -3679 381
rect -3617 347 -3583 381
rect -3521 347 -3487 381
rect -3425 347 -3391 381
rect -3329 347 -3295 381
rect -3233 347 -3199 381
rect -3137 347 -3103 381
rect -3041 347 -3007 381
rect -2945 347 -2911 381
rect -2849 347 -2815 381
rect -2753 347 -2719 381
rect -2657 347 -2623 381
rect -2561 347 -2527 381
rect -2465 347 -2431 381
rect -2369 347 -2335 381
rect -2273 347 -2239 381
rect -2177 347 -2143 381
rect -2081 347 -2047 381
rect -1985 347 -1951 381
rect -1889 347 -1855 381
rect -1793 347 -1759 381
rect -1697 347 -1663 381
rect -1601 347 -1567 381
rect -1505 347 -1471 381
rect -1409 347 -1375 381
rect -1313 347 -1279 381
rect -1217 347 -1183 381
rect -1121 347 -1087 381
rect -1025 347 -991 381
rect -929 347 -895 381
rect -833 347 -799 381
rect -737 347 -703 381
rect -641 347 -607 381
rect -545 347 -511 381
rect -449 347 -415 381
rect -353 347 -319 381
rect -257 347 -223 381
rect -161 347 -127 381
rect -65 347 -31 381
rect 31 347 65 381
rect 127 347 161 381
rect 223 347 257 381
rect 319 347 353 381
rect 415 347 449 381
rect 511 347 545 381
rect 607 347 641 381
rect 703 347 737 381
rect 799 347 833 381
rect 895 347 929 381
rect 991 347 1025 381
rect 1087 347 1121 381
rect 1183 347 1217 381
rect 1279 347 1313 381
rect 1375 347 1409 381
rect 1471 347 1505 381
rect 1567 347 1601 381
rect 1663 347 1697 381
rect 1759 347 1793 381
rect 1855 347 1889 381
rect 1951 347 1985 381
rect 2047 347 2081 381
rect 2143 347 2177 381
rect 2239 347 2273 381
rect 2335 347 2369 381
rect 2431 347 2465 381
rect 2527 347 2561 381
rect 2623 347 2657 381
rect 2719 347 2753 381
rect 2815 347 2849 381
rect 2911 347 2945 381
rect 3007 347 3041 381
rect 3103 347 3137 381
rect 3199 347 3233 381
rect 3295 347 3329 381
rect 3391 347 3425 381
rect 3487 347 3521 381
rect 3583 347 3617 381
rect 3679 347 3713 381
rect 3775 347 3809 381
rect 3871 347 3905 381
rect 3967 347 4001 381
rect 4063 347 4097 381
rect 4159 347 4193 381
rect 4255 347 4289 381
rect 4351 347 4385 381
rect 4447 347 4481 381
rect 4543 347 4577 381
rect 4639 347 4673 381
rect 4735 347 4769 381
rect 4831 347 4865 381
rect 4927 347 4961 381
rect 5023 347 5057 381
rect 5119 347 5153 381
rect 5215 347 5249 381
rect 5311 347 5345 381
rect 5407 347 5441 381
rect 5503 347 5537 381
rect 5599 347 5633 381
rect 5695 347 5729 381
rect -5777 -288 -5743 288
rect -5681 -288 -5647 288
rect -5585 -288 -5551 288
rect -5489 -288 -5455 288
rect -5393 -288 -5359 288
rect -5297 -288 -5263 288
rect -5201 -288 -5167 288
rect -5105 -288 -5071 288
rect -5009 -288 -4975 288
rect -4913 -288 -4879 288
rect -4817 -288 -4783 288
rect -4721 -288 -4687 288
rect -4625 -288 -4591 288
rect -4529 -288 -4495 288
rect -4433 -288 -4399 288
rect -4337 -288 -4303 288
rect -4241 -288 -4207 288
rect -4145 -288 -4111 288
rect -4049 -288 -4015 288
rect -3953 -288 -3919 288
rect -3857 -288 -3823 288
rect -3761 -288 -3727 288
rect -3665 -288 -3631 288
rect -3569 -288 -3535 288
rect -3473 -288 -3439 288
rect -3377 -288 -3343 288
rect -3281 -288 -3247 288
rect -3185 -288 -3151 288
rect -3089 -288 -3055 288
rect -2993 -288 -2959 288
rect -2897 -288 -2863 288
rect -2801 -288 -2767 288
rect -2705 -288 -2671 288
rect -2609 -288 -2575 288
rect -2513 -288 -2479 288
rect -2417 -288 -2383 288
rect -2321 -288 -2287 288
rect -2225 -288 -2191 288
rect -2129 -288 -2095 288
rect -2033 -288 -1999 288
rect -1937 -288 -1903 288
rect -1841 -288 -1807 288
rect -1745 -288 -1711 288
rect -1649 -288 -1615 288
rect -1553 -288 -1519 288
rect -1457 -288 -1423 288
rect -1361 -288 -1327 288
rect -1265 -288 -1231 288
rect -1169 -288 -1135 288
rect -1073 -288 -1039 288
rect -977 -288 -943 288
rect -881 -288 -847 288
rect -785 -288 -751 288
rect -689 -288 -655 288
rect -593 -288 -559 288
rect -497 -288 -463 288
rect -401 -288 -367 288
rect -305 -288 -271 288
rect -209 -288 -175 288
rect -113 -288 -79 288
rect -17 -288 17 288
rect 79 -288 113 288
rect 175 -288 209 288
rect 271 -288 305 288
rect 367 -288 401 288
rect 463 -288 497 288
rect 559 -288 593 288
rect 655 -288 689 288
rect 751 -288 785 288
rect 847 -288 881 288
rect 943 -288 977 288
rect 1039 -288 1073 288
rect 1135 -288 1169 288
rect 1231 -288 1265 288
rect 1327 -288 1361 288
rect 1423 -288 1457 288
rect 1519 -288 1553 288
rect 1615 -288 1649 288
rect 1711 -288 1745 288
rect 1807 -288 1841 288
rect 1903 -288 1937 288
rect 1999 -288 2033 288
rect 2095 -288 2129 288
rect 2191 -288 2225 288
rect 2287 -288 2321 288
rect 2383 -288 2417 288
rect 2479 -288 2513 288
rect 2575 -288 2609 288
rect 2671 -288 2705 288
rect 2767 -288 2801 288
rect 2863 -288 2897 288
rect 2959 -288 2993 288
rect 3055 -288 3089 288
rect 3151 -288 3185 288
rect 3247 -288 3281 288
rect 3343 -288 3377 288
rect 3439 -288 3473 288
rect 3535 -288 3569 288
rect 3631 -288 3665 288
rect 3727 -288 3761 288
rect 3823 -288 3857 288
rect 3919 -288 3953 288
rect 4015 -288 4049 288
rect 4111 -288 4145 288
rect 4207 -288 4241 288
rect 4303 -288 4337 288
rect 4399 -288 4433 288
rect 4495 -288 4529 288
rect 4591 -288 4625 288
rect 4687 -288 4721 288
rect 4783 -288 4817 288
rect 4879 -288 4913 288
rect 4975 -288 5009 288
rect 5071 -288 5105 288
rect 5167 -288 5201 288
rect 5263 -288 5297 288
rect 5359 -288 5393 288
rect 5455 -288 5489 288
rect 5551 -288 5585 288
rect 5647 -288 5681 288
rect 5743 -288 5777 288
rect -5729 -381 -5695 -347
rect -5633 -381 -5599 -347
rect -5537 -381 -5503 -347
rect -5441 -381 -5407 -347
rect -5345 -381 -5311 -347
rect -5249 -381 -5215 -347
rect -5153 -381 -5119 -347
rect -5057 -381 -5023 -347
rect -4961 -381 -4927 -347
rect -4865 -381 -4831 -347
rect -4769 -381 -4735 -347
rect -4673 -381 -4639 -347
rect -4577 -381 -4543 -347
rect -4481 -381 -4447 -347
rect -4385 -381 -4351 -347
rect -4289 -381 -4255 -347
rect -4193 -381 -4159 -347
rect -4097 -381 -4063 -347
rect -4001 -381 -3967 -347
rect -3905 -381 -3871 -347
rect -3809 -381 -3775 -347
rect -3713 -381 -3679 -347
rect -3617 -381 -3583 -347
rect -3521 -381 -3487 -347
rect -3425 -381 -3391 -347
rect -3329 -381 -3295 -347
rect -3233 -381 -3199 -347
rect -3137 -381 -3103 -347
rect -3041 -381 -3007 -347
rect -2945 -381 -2911 -347
rect -2849 -381 -2815 -347
rect -2753 -381 -2719 -347
rect -2657 -381 -2623 -347
rect -2561 -381 -2527 -347
rect -2465 -381 -2431 -347
rect -2369 -381 -2335 -347
rect -2273 -381 -2239 -347
rect -2177 -381 -2143 -347
rect -2081 -381 -2047 -347
rect -1985 -381 -1951 -347
rect -1889 -381 -1855 -347
rect -1793 -381 -1759 -347
rect -1697 -381 -1663 -347
rect -1601 -381 -1567 -347
rect -1505 -381 -1471 -347
rect -1409 -381 -1375 -347
rect -1313 -381 -1279 -347
rect -1217 -381 -1183 -347
rect -1121 -381 -1087 -347
rect -1025 -381 -991 -347
rect -929 -381 -895 -347
rect -833 -381 -799 -347
rect -737 -381 -703 -347
rect -641 -381 -607 -347
rect -545 -381 -511 -347
rect -449 -381 -415 -347
rect -353 -381 -319 -347
rect -257 -381 -223 -347
rect -161 -381 -127 -347
rect -65 -381 -31 -347
rect 31 -381 65 -347
rect 127 -381 161 -347
rect 223 -381 257 -347
rect 319 -381 353 -347
rect 415 -381 449 -347
rect 511 -381 545 -347
rect 607 -381 641 -347
rect 703 -381 737 -347
rect 799 -381 833 -347
rect 895 -381 929 -347
rect 991 -381 1025 -347
rect 1087 -381 1121 -347
rect 1183 -381 1217 -347
rect 1279 -381 1313 -347
rect 1375 -381 1409 -347
rect 1471 -381 1505 -347
rect 1567 -381 1601 -347
rect 1663 -381 1697 -347
rect 1759 -381 1793 -347
rect 1855 -381 1889 -347
rect 1951 -381 1985 -347
rect 2047 -381 2081 -347
rect 2143 -381 2177 -347
rect 2239 -381 2273 -347
rect 2335 -381 2369 -347
rect 2431 -381 2465 -347
rect 2527 -381 2561 -347
rect 2623 -381 2657 -347
rect 2719 -381 2753 -347
rect 2815 -381 2849 -347
rect 2911 -381 2945 -347
rect 3007 -381 3041 -347
rect 3103 -381 3137 -347
rect 3199 -381 3233 -347
rect 3295 -381 3329 -347
rect 3391 -381 3425 -347
rect 3487 -381 3521 -347
rect 3583 -381 3617 -347
rect 3679 -381 3713 -347
rect 3775 -381 3809 -347
rect 3871 -381 3905 -347
rect 3967 -381 4001 -347
rect 4063 -381 4097 -347
rect 4159 -381 4193 -347
rect 4255 -381 4289 -347
rect 4351 -381 4385 -347
rect 4447 -381 4481 -347
rect 4543 -381 4577 -347
rect 4639 -381 4673 -347
rect 4735 -381 4769 -347
rect 4831 -381 4865 -347
rect 4927 -381 4961 -347
rect 5023 -381 5057 -347
rect 5119 -381 5153 -347
rect 5215 -381 5249 -347
rect 5311 -381 5345 -347
rect 5407 -381 5441 -347
rect 5503 -381 5537 -347
rect 5599 -381 5633 -347
rect 5695 -381 5729 -347
rect 5857 -387 5891 387
rect -5885 -483 -5795 -449
rect -5795 -483 5795 -449
<< metal1 >>
rect -5897 483 5897 489
rect -5897 449 -5885 483
rect 5795 449 5897 483
rect -5897 443 5897 449
rect 5851 387 5897 443
rect -5897 381 5741 387
rect -5897 347 -5729 381
rect -5695 347 -5633 381
rect -5599 347 -5537 381
rect -5503 347 -5441 381
rect -5407 347 -5345 381
rect -5311 347 -5249 381
rect -5215 347 -5153 381
rect -5119 347 -5057 381
rect -5023 347 -4961 381
rect -4927 347 -4865 381
rect -4831 347 -4769 381
rect -4735 347 -4673 381
rect -4639 347 -4577 381
rect -4543 347 -4481 381
rect -4447 347 -4385 381
rect -4351 347 -4289 381
rect -4255 347 -4193 381
rect -4159 347 -4097 381
rect -4063 347 -4001 381
rect -3967 347 -3905 381
rect -3871 347 -3809 381
rect -3775 347 -3713 381
rect -3679 347 -3617 381
rect -3583 347 -3521 381
rect -3487 347 -3425 381
rect -3391 347 -3329 381
rect -3295 347 -3233 381
rect -3199 347 -3137 381
rect -3103 347 -3041 381
rect -3007 347 -2945 381
rect -2911 347 -2849 381
rect -2815 347 -2753 381
rect -2719 347 -2657 381
rect -2623 347 -2561 381
rect -2527 347 -2465 381
rect -2431 347 -2369 381
rect -2335 347 -2273 381
rect -2239 347 -2177 381
rect -2143 347 -2081 381
rect -2047 347 -1985 381
rect -1951 347 -1889 381
rect -1855 347 -1793 381
rect -1759 347 -1697 381
rect -1663 347 -1601 381
rect -1567 347 -1505 381
rect -1471 347 -1409 381
rect -1375 347 -1313 381
rect -1279 347 -1217 381
rect -1183 347 -1121 381
rect -1087 347 -1025 381
rect -991 347 -929 381
rect -895 347 -833 381
rect -799 347 -737 381
rect -703 347 -641 381
rect -607 347 -545 381
rect -511 347 -449 381
rect -415 347 -353 381
rect -319 347 -257 381
rect -223 347 -161 381
rect -127 347 -65 381
rect -31 347 31 381
rect 65 347 127 381
rect 161 347 223 381
rect 257 347 319 381
rect 353 347 415 381
rect 449 347 511 381
rect 545 347 607 381
rect 641 347 703 381
rect 737 347 799 381
rect 833 347 895 381
rect 929 347 991 381
rect 1025 347 1087 381
rect 1121 347 1183 381
rect 1217 347 1279 381
rect 1313 347 1375 381
rect 1409 347 1471 381
rect 1505 347 1567 381
rect 1601 347 1663 381
rect 1697 347 1759 381
rect 1793 347 1855 381
rect 1889 347 1951 381
rect 1985 347 2047 381
rect 2081 347 2143 381
rect 2177 347 2239 381
rect 2273 347 2335 381
rect 2369 347 2431 381
rect 2465 347 2527 381
rect 2561 347 2623 381
rect 2657 347 2719 381
rect 2753 347 2815 381
rect 2849 347 2911 381
rect 2945 347 3007 381
rect 3041 347 3103 381
rect 3137 347 3199 381
rect 3233 347 3295 381
rect 3329 347 3391 381
rect 3425 347 3487 381
rect 3521 347 3583 381
rect 3617 347 3679 381
rect 3713 347 3775 381
rect 3809 347 3871 381
rect 3905 347 3967 381
rect 4001 347 4063 381
rect 4097 347 4159 381
rect 4193 347 4255 381
rect 4289 347 4351 381
rect 4385 347 4447 381
rect 4481 347 4543 381
rect 4577 347 4639 381
rect 4673 347 4735 381
rect 4769 347 4831 381
rect 4865 347 4927 381
rect 4961 347 5023 381
rect 5057 347 5119 381
rect 5153 347 5215 381
rect 5249 347 5311 381
rect 5345 347 5407 381
rect 5441 347 5503 381
rect 5537 347 5599 381
rect 5633 347 5695 381
rect 5729 347 5741 381
rect -5897 341 5741 347
rect -5897 -341 -5851 341
rect -5786 288 -5734 300
rect -5786 -26 -5777 288
rect -5743 -26 -5734 288
rect -5786 -300 -5734 -294
rect -5690 294 -5638 300
rect -5690 -288 -5681 26
rect -5647 -288 -5638 26
rect -5690 -300 -5638 -288
rect -5594 288 -5542 300
rect -5594 -26 -5585 288
rect -5551 -26 -5542 288
rect -5594 -300 -5542 -294
rect -5498 294 -5446 300
rect -5498 -288 -5489 26
rect -5455 -288 -5446 26
rect -5498 -300 -5446 -288
rect -5402 288 -5350 300
rect -5402 -26 -5393 288
rect -5359 -26 -5350 288
rect -5402 -300 -5350 -294
rect -5306 294 -5254 300
rect -5306 -288 -5297 26
rect -5263 -288 -5254 26
rect -5306 -300 -5254 -288
rect -5210 288 -5158 300
rect -5210 -26 -5201 288
rect -5167 -26 -5158 288
rect -5210 -300 -5158 -294
rect -5114 294 -5062 300
rect -5114 -288 -5105 26
rect -5071 -288 -5062 26
rect -5114 -300 -5062 -288
rect -5018 288 -4966 300
rect -5018 -26 -5009 288
rect -4975 -26 -4966 288
rect -5018 -300 -4966 -294
rect -4922 294 -4870 300
rect -4922 -288 -4913 26
rect -4879 -288 -4870 26
rect -4922 -300 -4870 -288
rect -4826 288 -4774 300
rect -4826 -26 -4817 288
rect -4783 -26 -4774 288
rect -4826 -300 -4774 -294
rect -4730 294 -4678 300
rect -4730 -288 -4721 26
rect -4687 -288 -4678 26
rect -4730 -300 -4678 -288
rect -4634 288 -4582 300
rect -4634 -26 -4625 288
rect -4591 -26 -4582 288
rect -4634 -300 -4582 -294
rect -4538 294 -4486 300
rect -4538 -288 -4529 26
rect -4495 -288 -4486 26
rect -4538 -300 -4486 -288
rect -4442 288 -4390 300
rect -4442 -26 -4433 288
rect -4399 -26 -4390 288
rect -4442 -300 -4390 -294
rect -4346 294 -4294 300
rect -4346 -288 -4337 26
rect -4303 -288 -4294 26
rect -4346 -300 -4294 -288
rect -4250 288 -4198 300
rect -4250 -26 -4241 288
rect -4207 -26 -4198 288
rect -4250 -300 -4198 -294
rect -4154 294 -4102 300
rect -4154 -288 -4145 26
rect -4111 -288 -4102 26
rect -4154 -300 -4102 -288
rect -4058 288 -4006 300
rect -4058 -26 -4049 288
rect -4015 -26 -4006 288
rect -4058 -300 -4006 -294
rect -3962 294 -3910 300
rect -3962 -288 -3953 26
rect -3919 -288 -3910 26
rect -3962 -300 -3910 -288
rect -3866 288 -3814 300
rect -3866 -26 -3857 288
rect -3823 -26 -3814 288
rect -3866 -300 -3814 -294
rect -3770 294 -3718 300
rect -3770 -288 -3761 26
rect -3727 -288 -3718 26
rect -3770 -300 -3718 -288
rect -3674 288 -3622 300
rect -3674 -26 -3665 288
rect -3631 -26 -3622 288
rect -3674 -300 -3622 -294
rect -3578 294 -3526 300
rect -3578 -288 -3569 26
rect -3535 -288 -3526 26
rect -3578 -300 -3526 -288
rect -3482 288 -3430 300
rect -3482 -26 -3473 288
rect -3439 -26 -3430 288
rect -3482 -300 -3430 -294
rect -3386 294 -3334 300
rect -3386 -288 -3377 26
rect -3343 -288 -3334 26
rect -3386 -300 -3334 -288
rect -3290 288 -3238 300
rect -3290 -26 -3281 288
rect -3247 -26 -3238 288
rect -3290 -300 -3238 -294
rect -3194 294 -3142 300
rect -3194 -288 -3185 26
rect -3151 -288 -3142 26
rect -3194 -300 -3142 -288
rect -3098 288 -3046 300
rect -3098 -26 -3089 288
rect -3055 -26 -3046 288
rect -3098 -300 -3046 -294
rect -3002 294 -2950 300
rect -3002 -288 -2993 26
rect -2959 -288 -2950 26
rect -3002 -300 -2950 -288
rect -2906 288 -2854 300
rect -2906 -26 -2897 288
rect -2863 -26 -2854 288
rect -2906 -300 -2854 -294
rect -2810 294 -2758 300
rect -2810 -288 -2801 26
rect -2767 -288 -2758 26
rect -2810 -300 -2758 -288
rect -2714 288 -2662 300
rect -2714 -26 -2705 288
rect -2671 -26 -2662 288
rect -2714 -300 -2662 -294
rect -2618 294 -2566 300
rect -2618 -288 -2609 26
rect -2575 -288 -2566 26
rect -2618 -300 -2566 -288
rect -2522 288 -2470 300
rect -2522 -26 -2513 288
rect -2479 -26 -2470 288
rect -2522 -300 -2470 -294
rect -2426 294 -2374 300
rect -2426 -288 -2417 26
rect -2383 -288 -2374 26
rect -2426 -300 -2374 -288
rect -2330 288 -2278 300
rect -2330 -26 -2321 288
rect -2287 -26 -2278 288
rect -2330 -300 -2278 -294
rect -2234 294 -2182 300
rect -2234 -288 -2225 26
rect -2191 -288 -2182 26
rect -2234 -300 -2182 -288
rect -2138 288 -2086 300
rect -2138 -26 -2129 288
rect -2095 -26 -2086 288
rect -2138 -300 -2086 -294
rect -2042 294 -1990 300
rect -2042 -288 -2033 26
rect -1999 -288 -1990 26
rect -2042 -300 -1990 -288
rect -1946 288 -1894 300
rect -1946 -26 -1937 288
rect -1903 -26 -1894 288
rect -1946 -300 -1894 -294
rect -1850 294 -1798 300
rect -1850 -288 -1841 26
rect -1807 -288 -1798 26
rect -1850 -300 -1798 -288
rect -1754 288 -1702 300
rect -1754 -26 -1745 288
rect -1711 -26 -1702 288
rect -1754 -300 -1702 -294
rect -1658 294 -1606 300
rect -1658 -288 -1649 26
rect -1615 -288 -1606 26
rect -1658 -300 -1606 -288
rect -1562 288 -1510 300
rect -1562 -26 -1553 288
rect -1519 -26 -1510 288
rect -1562 -300 -1510 -294
rect -1466 294 -1414 300
rect -1466 -288 -1457 26
rect -1423 -288 -1414 26
rect -1466 -300 -1414 -288
rect -1370 288 -1318 300
rect -1370 -26 -1361 288
rect -1327 -26 -1318 288
rect -1370 -300 -1318 -294
rect -1274 294 -1222 300
rect -1274 -288 -1265 26
rect -1231 -288 -1222 26
rect -1274 -300 -1222 -288
rect -1178 288 -1126 300
rect -1178 -26 -1169 288
rect -1135 -26 -1126 288
rect -1178 -300 -1126 -294
rect -1082 294 -1030 300
rect -1082 -288 -1073 26
rect -1039 -288 -1030 26
rect -1082 -300 -1030 -288
rect -986 288 -934 300
rect -986 -26 -977 288
rect -943 -26 -934 288
rect -986 -300 -934 -294
rect -890 294 -838 300
rect -890 -288 -881 26
rect -847 -288 -838 26
rect -890 -300 -838 -288
rect -794 288 -742 300
rect -794 -26 -785 288
rect -751 -26 -742 288
rect -794 -300 -742 -294
rect -698 294 -646 300
rect -698 -288 -689 26
rect -655 -288 -646 26
rect -698 -300 -646 -288
rect -602 288 -550 300
rect -602 -26 -593 288
rect -559 -26 -550 288
rect -602 -300 -550 -294
rect -506 294 -454 300
rect -506 -288 -497 26
rect -463 -288 -454 26
rect -506 -300 -454 -288
rect -410 288 -358 300
rect -410 -26 -401 288
rect -367 -26 -358 288
rect -410 -300 -358 -294
rect -314 294 -262 300
rect -314 -288 -305 26
rect -271 -288 -262 26
rect -314 -300 -262 -288
rect -218 288 -166 300
rect -218 -26 -209 288
rect -175 -26 -166 288
rect -218 -300 -166 -294
rect -122 294 -70 300
rect -122 -288 -113 26
rect -79 -288 -70 26
rect -122 -300 -70 -288
rect -26 288 26 300
rect -26 -26 -17 288
rect 17 -26 26 288
rect -26 -300 26 -294
rect 70 294 122 300
rect 70 -288 79 26
rect 113 -288 122 26
rect 70 -300 122 -288
rect 166 288 218 300
rect 166 -26 175 288
rect 209 -26 218 288
rect 166 -300 218 -294
rect 262 294 314 300
rect 262 -288 271 26
rect 305 -288 314 26
rect 262 -300 314 -288
rect 358 288 410 300
rect 358 -26 367 288
rect 401 -26 410 288
rect 358 -300 410 -294
rect 454 294 506 300
rect 454 -288 463 26
rect 497 -288 506 26
rect 454 -300 506 -288
rect 550 288 602 300
rect 550 -26 559 288
rect 593 -26 602 288
rect 550 -300 602 -294
rect 646 294 698 300
rect 646 -288 655 26
rect 689 -288 698 26
rect 646 -300 698 -288
rect 742 288 794 300
rect 742 -26 751 288
rect 785 -26 794 288
rect 742 -300 794 -294
rect 838 294 890 300
rect 838 -288 847 26
rect 881 -288 890 26
rect 838 -300 890 -288
rect 934 288 986 300
rect 934 -26 943 288
rect 977 -26 986 288
rect 934 -300 986 -294
rect 1030 294 1082 300
rect 1030 -288 1039 26
rect 1073 -288 1082 26
rect 1030 -300 1082 -288
rect 1126 288 1178 300
rect 1126 -26 1135 288
rect 1169 -26 1178 288
rect 1126 -300 1178 -294
rect 1222 294 1274 300
rect 1222 -288 1231 26
rect 1265 -288 1274 26
rect 1222 -300 1274 -288
rect 1318 288 1370 300
rect 1318 -26 1327 288
rect 1361 -26 1370 288
rect 1318 -300 1370 -294
rect 1414 294 1466 300
rect 1414 -288 1423 26
rect 1457 -288 1466 26
rect 1414 -300 1466 -288
rect 1510 288 1562 300
rect 1510 -26 1519 288
rect 1553 -26 1562 288
rect 1510 -300 1562 -294
rect 1606 294 1658 300
rect 1606 -288 1615 26
rect 1649 -288 1658 26
rect 1606 -300 1658 -288
rect 1702 288 1754 300
rect 1702 -26 1711 288
rect 1745 -26 1754 288
rect 1702 -300 1754 -294
rect 1798 294 1850 300
rect 1798 -288 1807 26
rect 1841 -288 1850 26
rect 1798 -300 1850 -288
rect 1894 288 1946 300
rect 1894 -26 1903 288
rect 1937 -26 1946 288
rect 1894 -300 1946 -294
rect 1990 294 2042 300
rect 1990 -288 1999 26
rect 2033 -288 2042 26
rect 1990 -300 2042 -288
rect 2086 288 2138 300
rect 2086 -26 2095 288
rect 2129 -26 2138 288
rect 2086 -300 2138 -294
rect 2182 294 2234 300
rect 2182 -288 2191 26
rect 2225 -288 2234 26
rect 2182 -300 2234 -288
rect 2278 288 2330 300
rect 2278 -26 2287 288
rect 2321 -26 2330 288
rect 2278 -300 2330 -294
rect 2374 294 2426 300
rect 2374 -288 2383 26
rect 2417 -288 2426 26
rect 2374 -300 2426 -288
rect 2470 288 2522 300
rect 2470 -26 2479 288
rect 2513 -26 2522 288
rect 2470 -300 2522 -294
rect 2566 294 2618 300
rect 2566 -288 2575 26
rect 2609 -288 2618 26
rect 2566 -300 2618 -288
rect 2662 288 2714 300
rect 2662 -26 2671 288
rect 2705 -26 2714 288
rect 2662 -300 2714 -294
rect 2758 294 2810 300
rect 2758 -288 2767 26
rect 2801 -288 2810 26
rect 2758 -300 2810 -288
rect 2854 288 2906 300
rect 2854 -26 2863 288
rect 2897 -26 2906 288
rect 2854 -300 2906 -294
rect 2950 294 3002 300
rect 2950 -288 2959 26
rect 2993 -288 3002 26
rect 2950 -300 3002 -288
rect 3046 288 3098 300
rect 3046 -26 3055 288
rect 3089 -26 3098 288
rect 3046 -300 3098 -294
rect 3142 294 3194 300
rect 3142 -288 3151 26
rect 3185 -288 3194 26
rect 3142 -300 3194 -288
rect 3238 288 3290 300
rect 3238 -26 3247 288
rect 3281 -26 3290 288
rect 3238 -300 3290 -294
rect 3334 294 3386 300
rect 3334 -288 3343 26
rect 3377 -288 3386 26
rect 3334 -300 3386 -288
rect 3430 288 3482 300
rect 3430 -26 3439 288
rect 3473 -26 3482 288
rect 3430 -300 3482 -294
rect 3526 294 3578 300
rect 3526 -288 3535 26
rect 3569 -288 3578 26
rect 3526 -300 3578 -288
rect 3622 288 3674 300
rect 3622 -26 3631 288
rect 3665 -26 3674 288
rect 3622 -300 3674 -294
rect 3718 294 3770 300
rect 3718 -288 3727 26
rect 3761 -288 3770 26
rect 3718 -300 3770 -288
rect 3814 288 3866 300
rect 3814 -26 3823 288
rect 3857 -26 3866 288
rect 3814 -300 3866 -294
rect 3910 294 3962 300
rect 3910 -288 3919 26
rect 3953 -288 3962 26
rect 3910 -300 3962 -288
rect 4006 288 4058 300
rect 4006 -26 4015 288
rect 4049 -26 4058 288
rect 4006 -300 4058 -294
rect 4102 294 4154 300
rect 4102 -288 4111 26
rect 4145 -288 4154 26
rect 4102 -300 4154 -288
rect 4198 288 4250 300
rect 4198 -26 4207 288
rect 4241 -26 4250 288
rect 4198 -300 4250 -294
rect 4294 294 4346 300
rect 4294 -288 4303 26
rect 4337 -288 4346 26
rect 4294 -300 4346 -288
rect 4390 288 4442 300
rect 4390 -26 4399 288
rect 4433 -26 4442 288
rect 4390 -300 4442 -294
rect 4486 294 4538 300
rect 4486 -288 4495 26
rect 4529 -288 4538 26
rect 4486 -300 4538 -288
rect 4582 288 4634 300
rect 4582 -26 4591 288
rect 4625 -26 4634 288
rect 4582 -300 4634 -294
rect 4678 294 4730 300
rect 4678 -288 4687 26
rect 4721 -288 4730 26
rect 4678 -300 4730 -288
rect 4774 288 4826 300
rect 4774 -26 4783 288
rect 4817 -26 4826 288
rect 4774 -300 4826 -294
rect 4870 294 4922 300
rect 4870 -288 4879 26
rect 4913 -288 4922 26
rect 4870 -300 4922 -288
rect 4966 288 5018 300
rect 4966 -26 4975 288
rect 5009 -26 5018 288
rect 4966 -300 5018 -294
rect 5062 294 5114 300
rect 5062 -288 5071 26
rect 5105 -288 5114 26
rect 5062 -300 5114 -288
rect 5158 288 5210 300
rect 5158 -26 5167 288
rect 5201 -26 5210 288
rect 5158 -300 5210 -294
rect 5254 294 5306 300
rect 5254 -288 5263 26
rect 5297 -288 5306 26
rect 5254 -300 5306 -288
rect 5350 288 5402 300
rect 5350 -26 5359 288
rect 5393 -26 5402 288
rect 5350 -300 5402 -294
rect 5446 294 5498 300
rect 5446 -288 5455 26
rect 5489 -288 5498 26
rect 5446 -300 5498 -288
rect 5542 288 5594 300
rect 5542 -26 5551 288
rect 5585 -26 5594 288
rect 5542 -300 5594 -294
rect 5638 294 5690 300
rect 5638 -288 5647 26
rect 5681 -288 5690 26
rect 5638 -300 5690 -288
rect 5734 288 5786 300
rect 5734 -26 5743 288
rect 5777 -26 5786 288
rect 5734 -300 5786 -294
rect -5897 -347 5741 -341
rect -5897 -381 -5729 -347
rect -5695 -381 -5633 -347
rect -5599 -381 -5537 -347
rect -5503 -381 -5441 -347
rect -5407 -381 -5345 -347
rect -5311 -381 -5249 -347
rect -5215 -381 -5153 -347
rect -5119 -381 -5057 -347
rect -5023 -381 -4961 -347
rect -4927 -381 -4865 -347
rect -4831 -381 -4769 -347
rect -4735 -381 -4673 -347
rect -4639 -381 -4577 -347
rect -4543 -381 -4481 -347
rect -4447 -381 -4385 -347
rect -4351 -381 -4289 -347
rect -4255 -381 -4193 -347
rect -4159 -381 -4097 -347
rect -4063 -381 -4001 -347
rect -3967 -381 -3905 -347
rect -3871 -381 -3809 -347
rect -3775 -381 -3713 -347
rect -3679 -381 -3617 -347
rect -3583 -381 -3521 -347
rect -3487 -381 -3425 -347
rect -3391 -381 -3329 -347
rect -3295 -381 -3233 -347
rect -3199 -381 -3137 -347
rect -3103 -381 -3041 -347
rect -3007 -381 -2945 -347
rect -2911 -381 -2849 -347
rect -2815 -381 -2753 -347
rect -2719 -381 -2657 -347
rect -2623 -381 -2561 -347
rect -2527 -381 -2465 -347
rect -2431 -381 -2369 -347
rect -2335 -381 -2273 -347
rect -2239 -381 -2177 -347
rect -2143 -381 -2081 -347
rect -2047 -381 -1985 -347
rect -1951 -381 -1889 -347
rect -1855 -381 -1793 -347
rect -1759 -381 -1697 -347
rect -1663 -381 -1601 -347
rect -1567 -381 -1505 -347
rect -1471 -381 -1409 -347
rect -1375 -381 -1313 -347
rect -1279 -381 -1217 -347
rect -1183 -381 -1121 -347
rect -1087 -381 -1025 -347
rect -991 -381 -929 -347
rect -895 -381 -833 -347
rect -799 -381 -737 -347
rect -703 -381 -641 -347
rect -607 -381 -545 -347
rect -511 -381 -449 -347
rect -415 -381 -353 -347
rect -319 -381 -257 -347
rect -223 -381 -161 -347
rect -127 -381 -65 -347
rect -31 -381 31 -347
rect 65 -381 127 -347
rect 161 -381 223 -347
rect 257 -381 319 -347
rect 353 -381 415 -347
rect 449 -381 511 -347
rect 545 -381 607 -347
rect 641 -381 703 -347
rect 737 -381 799 -347
rect 833 -381 895 -347
rect 929 -381 991 -347
rect 1025 -381 1087 -347
rect 1121 -381 1183 -347
rect 1217 -381 1279 -347
rect 1313 -381 1375 -347
rect 1409 -381 1471 -347
rect 1505 -381 1567 -347
rect 1601 -381 1663 -347
rect 1697 -381 1759 -347
rect 1793 -381 1855 -347
rect 1889 -381 1951 -347
rect 1985 -381 2047 -347
rect 2081 -381 2143 -347
rect 2177 -381 2239 -347
rect 2273 -381 2335 -347
rect 2369 -381 2431 -347
rect 2465 -381 2527 -347
rect 2561 -381 2623 -347
rect 2657 -381 2719 -347
rect 2753 -381 2815 -347
rect 2849 -381 2911 -347
rect 2945 -381 3007 -347
rect 3041 -381 3103 -347
rect 3137 -381 3199 -347
rect 3233 -381 3295 -347
rect 3329 -381 3391 -347
rect 3425 -381 3487 -347
rect 3521 -381 3583 -347
rect 3617 -381 3679 -347
rect 3713 -381 3775 -347
rect 3809 -381 3871 -347
rect 3905 -381 3967 -347
rect 4001 -381 4063 -347
rect 4097 -381 4159 -347
rect 4193 -381 4255 -347
rect 4289 -381 4351 -347
rect 4385 -381 4447 -347
rect 4481 -381 4543 -347
rect 4577 -381 4639 -347
rect 4673 -381 4735 -347
rect 4769 -381 4831 -347
rect 4865 -381 4927 -347
rect 4961 -381 5023 -347
rect 5057 -381 5119 -347
rect 5153 -381 5215 -347
rect 5249 -381 5311 -347
rect 5345 -381 5407 -347
rect 5441 -381 5503 -347
rect 5537 -381 5599 -347
rect 5633 -381 5695 -347
rect 5729 -381 5741 -347
rect -5897 -387 5741 -381
rect 5851 -387 5857 387
rect 5891 -387 5897 387
rect 5851 -443 5897 -387
rect -5897 -449 5897 -443
rect -5897 -483 -5885 -449
rect 5795 -483 5897 -449
rect -5897 -489 5897 -483
<< via1 >>
rect -5786 -288 -5777 -26
rect -5777 -288 -5743 -26
rect -5743 -288 -5734 -26
rect -5786 -294 -5734 -288
rect -5690 288 -5638 294
rect -5690 26 -5681 288
rect -5681 26 -5647 288
rect -5647 26 -5638 288
rect -5594 -288 -5585 -26
rect -5585 -288 -5551 -26
rect -5551 -288 -5542 -26
rect -5594 -294 -5542 -288
rect -5498 288 -5446 294
rect -5498 26 -5489 288
rect -5489 26 -5455 288
rect -5455 26 -5446 288
rect -5402 -288 -5393 -26
rect -5393 -288 -5359 -26
rect -5359 -288 -5350 -26
rect -5402 -294 -5350 -288
rect -5306 288 -5254 294
rect -5306 26 -5297 288
rect -5297 26 -5263 288
rect -5263 26 -5254 288
rect -5210 -288 -5201 -26
rect -5201 -288 -5167 -26
rect -5167 -288 -5158 -26
rect -5210 -294 -5158 -288
rect -5114 288 -5062 294
rect -5114 26 -5105 288
rect -5105 26 -5071 288
rect -5071 26 -5062 288
rect -5018 -288 -5009 -26
rect -5009 -288 -4975 -26
rect -4975 -288 -4966 -26
rect -5018 -294 -4966 -288
rect -4922 288 -4870 294
rect -4922 26 -4913 288
rect -4913 26 -4879 288
rect -4879 26 -4870 288
rect -4826 -288 -4817 -26
rect -4817 -288 -4783 -26
rect -4783 -288 -4774 -26
rect -4826 -294 -4774 -288
rect -4730 288 -4678 294
rect -4730 26 -4721 288
rect -4721 26 -4687 288
rect -4687 26 -4678 288
rect -4634 -288 -4625 -26
rect -4625 -288 -4591 -26
rect -4591 -288 -4582 -26
rect -4634 -294 -4582 -288
rect -4538 288 -4486 294
rect -4538 26 -4529 288
rect -4529 26 -4495 288
rect -4495 26 -4486 288
rect -4442 -288 -4433 -26
rect -4433 -288 -4399 -26
rect -4399 -288 -4390 -26
rect -4442 -294 -4390 -288
rect -4346 288 -4294 294
rect -4346 26 -4337 288
rect -4337 26 -4303 288
rect -4303 26 -4294 288
rect -4250 -288 -4241 -26
rect -4241 -288 -4207 -26
rect -4207 -288 -4198 -26
rect -4250 -294 -4198 -288
rect -4154 288 -4102 294
rect -4154 26 -4145 288
rect -4145 26 -4111 288
rect -4111 26 -4102 288
rect -4058 -288 -4049 -26
rect -4049 -288 -4015 -26
rect -4015 -288 -4006 -26
rect -4058 -294 -4006 -288
rect -3962 288 -3910 294
rect -3962 26 -3953 288
rect -3953 26 -3919 288
rect -3919 26 -3910 288
rect -3866 -288 -3857 -26
rect -3857 -288 -3823 -26
rect -3823 -288 -3814 -26
rect -3866 -294 -3814 -288
rect -3770 288 -3718 294
rect -3770 26 -3761 288
rect -3761 26 -3727 288
rect -3727 26 -3718 288
rect -3674 -288 -3665 -26
rect -3665 -288 -3631 -26
rect -3631 -288 -3622 -26
rect -3674 -294 -3622 -288
rect -3578 288 -3526 294
rect -3578 26 -3569 288
rect -3569 26 -3535 288
rect -3535 26 -3526 288
rect -3482 -288 -3473 -26
rect -3473 -288 -3439 -26
rect -3439 -288 -3430 -26
rect -3482 -294 -3430 -288
rect -3386 288 -3334 294
rect -3386 26 -3377 288
rect -3377 26 -3343 288
rect -3343 26 -3334 288
rect -3290 -288 -3281 -26
rect -3281 -288 -3247 -26
rect -3247 -288 -3238 -26
rect -3290 -294 -3238 -288
rect -3194 288 -3142 294
rect -3194 26 -3185 288
rect -3185 26 -3151 288
rect -3151 26 -3142 288
rect -3098 -288 -3089 -26
rect -3089 -288 -3055 -26
rect -3055 -288 -3046 -26
rect -3098 -294 -3046 -288
rect -3002 288 -2950 294
rect -3002 26 -2993 288
rect -2993 26 -2959 288
rect -2959 26 -2950 288
rect -2906 -288 -2897 -26
rect -2897 -288 -2863 -26
rect -2863 -288 -2854 -26
rect -2906 -294 -2854 -288
rect -2810 288 -2758 294
rect -2810 26 -2801 288
rect -2801 26 -2767 288
rect -2767 26 -2758 288
rect -2714 -288 -2705 -26
rect -2705 -288 -2671 -26
rect -2671 -288 -2662 -26
rect -2714 -294 -2662 -288
rect -2618 288 -2566 294
rect -2618 26 -2609 288
rect -2609 26 -2575 288
rect -2575 26 -2566 288
rect -2522 -288 -2513 -26
rect -2513 -288 -2479 -26
rect -2479 -288 -2470 -26
rect -2522 -294 -2470 -288
rect -2426 288 -2374 294
rect -2426 26 -2417 288
rect -2417 26 -2383 288
rect -2383 26 -2374 288
rect -2330 -288 -2321 -26
rect -2321 -288 -2287 -26
rect -2287 -288 -2278 -26
rect -2330 -294 -2278 -288
rect -2234 288 -2182 294
rect -2234 26 -2225 288
rect -2225 26 -2191 288
rect -2191 26 -2182 288
rect -2138 -288 -2129 -26
rect -2129 -288 -2095 -26
rect -2095 -288 -2086 -26
rect -2138 -294 -2086 -288
rect -2042 288 -1990 294
rect -2042 26 -2033 288
rect -2033 26 -1999 288
rect -1999 26 -1990 288
rect -1946 -288 -1937 -26
rect -1937 -288 -1903 -26
rect -1903 -288 -1894 -26
rect -1946 -294 -1894 -288
rect -1850 288 -1798 294
rect -1850 26 -1841 288
rect -1841 26 -1807 288
rect -1807 26 -1798 288
rect -1754 -288 -1745 -26
rect -1745 -288 -1711 -26
rect -1711 -288 -1702 -26
rect -1754 -294 -1702 -288
rect -1658 288 -1606 294
rect -1658 26 -1649 288
rect -1649 26 -1615 288
rect -1615 26 -1606 288
rect -1562 -288 -1553 -26
rect -1553 -288 -1519 -26
rect -1519 -288 -1510 -26
rect -1562 -294 -1510 -288
rect -1466 288 -1414 294
rect -1466 26 -1457 288
rect -1457 26 -1423 288
rect -1423 26 -1414 288
rect -1370 -288 -1361 -26
rect -1361 -288 -1327 -26
rect -1327 -288 -1318 -26
rect -1370 -294 -1318 -288
rect -1274 288 -1222 294
rect -1274 26 -1265 288
rect -1265 26 -1231 288
rect -1231 26 -1222 288
rect -1178 -288 -1169 -26
rect -1169 -288 -1135 -26
rect -1135 -288 -1126 -26
rect -1178 -294 -1126 -288
rect -1082 288 -1030 294
rect -1082 26 -1073 288
rect -1073 26 -1039 288
rect -1039 26 -1030 288
rect -986 -288 -977 -26
rect -977 -288 -943 -26
rect -943 -288 -934 -26
rect -986 -294 -934 -288
rect -890 288 -838 294
rect -890 26 -881 288
rect -881 26 -847 288
rect -847 26 -838 288
rect -794 -288 -785 -26
rect -785 -288 -751 -26
rect -751 -288 -742 -26
rect -794 -294 -742 -288
rect -698 288 -646 294
rect -698 26 -689 288
rect -689 26 -655 288
rect -655 26 -646 288
rect -602 -288 -593 -26
rect -593 -288 -559 -26
rect -559 -288 -550 -26
rect -602 -294 -550 -288
rect -506 288 -454 294
rect -506 26 -497 288
rect -497 26 -463 288
rect -463 26 -454 288
rect -410 -288 -401 -26
rect -401 -288 -367 -26
rect -367 -288 -358 -26
rect -410 -294 -358 -288
rect -314 288 -262 294
rect -314 26 -305 288
rect -305 26 -271 288
rect -271 26 -262 288
rect -218 -288 -209 -26
rect -209 -288 -175 -26
rect -175 -288 -166 -26
rect -218 -294 -166 -288
rect -122 288 -70 294
rect -122 26 -113 288
rect -113 26 -79 288
rect -79 26 -70 288
rect -26 -288 -17 -26
rect -17 -288 17 -26
rect 17 -288 26 -26
rect -26 -294 26 -288
rect 70 288 122 294
rect 70 26 79 288
rect 79 26 113 288
rect 113 26 122 288
rect 166 -288 175 -26
rect 175 -288 209 -26
rect 209 -288 218 -26
rect 166 -294 218 -288
rect 262 288 314 294
rect 262 26 271 288
rect 271 26 305 288
rect 305 26 314 288
rect 358 -288 367 -26
rect 367 -288 401 -26
rect 401 -288 410 -26
rect 358 -294 410 -288
rect 454 288 506 294
rect 454 26 463 288
rect 463 26 497 288
rect 497 26 506 288
rect 550 -288 559 -26
rect 559 -288 593 -26
rect 593 -288 602 -26
rect 550 -294 602 -288
rect 646 288 698 294
rect 646 26 655 288
rect 655 26 689 288
rect 689 26 698 288
rect 742 -288 751 -26
rect 751 -288 785 -26
rect 785 -288 794 -26
rect 742 -294 794 -288
rect 838 288 890 294
rect 838 26 847 288
rect 847 26 881 288
rect 881 26 890 288
rect 934 -288 943 -26
rect 943 -288 977 -26
rect 977 -288 986 -26
rect 934 -294 986 -288
rect 1030 288 1082 294
rect 1030 26 1039 288
rect 1039 26 1073 288
rect 1073 26 1082 288
rect 1126 -288 1135 -26
rect 1135 -288 1169 -26
rect 1169 -288 1178 -26
rect 1126 -294 1178 -288
rect 1222 288 1274 294
rect 1222 26 1231 288
rect 1231 26 1265 288
rect 1265 26 1274 288
rect 1318 -288 1327 -26
rect 1327 -288 1361 -26
rect 1361 -288 1370 -26
rect 1318 -294 1370 -288
rect 1414 288 1466 294
rect 1414 26 1423 288
rect 1423 26 1457 288
rect 1457 26 1466 288
rect 1510 -288 1519 -26
rect 1519 -288 1553 -26
rect 1553 -288 1562 -26
rect 1510 -294 1562 -288
rect 1606 288 1658 294
rect 1606 26 1615 288
rect 1615 26 1649 288
rect 1649 26 1658 288
rect 1702 -288 1711 -26
rect 1711 -288 1745 -26
rect 1745 -288 1754 -26
rect 1702 -294 1754 -288
rect 1798 288 1850 294
rect 1798 26 1807 288
rect 1807 26 1841 288
rect 1841 26 1850 288
rect 1894 -288 1903 -26
rect 1903 -288 1937 -26
rect 1937 -288 1946 -26
rect 1894 -294 1946 -288
rect 1990 288 2042 294
rect 1990 26 1999 288
rect 1999 26 2033 288
rect 2033 26 2042 288
rect 2086 -288 2095 -26
rect 2095 -288 2129 -26
rect 2129 -288 2138 -26
rect 2086 -294 2138 -288
rect 2182 288 2234 294
rect 2182 26 2191 288
rect 2191 26 2225 288
rect 2225 26 2234 288
rect 2278 -288 2287 -26
rect 2287 -288 2321 -26
rect 2321 -288 2330 -26
rect 2278 -294 2330 -288
rect 2374 288 2426 294
rect 2374 26 2383 288
rect 2383 26 2417 288
rect 2417 26 2426 288
rect 2470 -288 2479 -26
rect 2479 -288 2513 -26
rect 2513 -288 2522 -26
rect 2470 -294 2522 -288
rect 2566 288 2618 294
rect 2566 26 2575 288
rect 2575 26 2609 288
rect 2609 26 2618 288
rect 2662 -288 2671 -26
rect 2671 -288 2705 -26
rect 2705 -288 2714 -26
rect 2662 -294 2714 -288
rect 2758 288 2810 294
rect 2758 26 2767 288
rect 2767 26 2801 288
rect 2801 26 2810 288
rect 2854 -288 2863 -26
rect 2863 -288 2897 -26
rect 2897 -288 2906 -26
rect 2854 -294 2906 -288
rect 2950 288 3002 294
rect 2950 26 2959 288
rect 2959 26 2993 288
rect 2993 26 3002 288
rect 3046 -288 3055 -26
rect 3055 -288 3089 -26
rect 3089 -288 3098 -26
rect 3046 -294 3098 -288
rect 3142 288 3194 294
rect 3142 26 3151 288
rect 3151 26 3185 288
rect 3185 26 3194 288
rect 3238 -288 3247 -26
rect 3247 -288 3281 -26
rect 3281 -288 3290 -26
rect 3238 -294 3290 -288
rect 3334 288 3386 294
rect 3334 26 3343 288
rect 3343 26 3377 288
rect 3377 26 3386 288
rect 3430 -288 3439 -26
rect 3439 -288 3473 -26
rect 3473 -288 3482 -26
rect 3430 -294 3482 -288
rect 3526 288 3578 294
rect 3526 26 3535 288
rect 3535 26 3569 288
rect 3569 26 3578 288
rect 3622 -288 3631 -26
rect 3631 -288 3665 -26
rect 3665 -288 3674 -26
rect 3622 -294 3674 -288
rect 3718 288 3770 294
rect 3718 26 3727 288
rect 3727 26 3761 288
rect 3761 26 3770 288
rect 3814 -288 3823 -26
rect 3823 -288 3857 -26
rect 3857 -288 3866 -26
rect 3814 -294 3866 -288
rect 3910 288 3962 294
rect 3910 26 3919 288
rect 3919 26 3953 288
rect 3953 26 3962 288
rect 4006 -288 4015 -26
rect 4015 -288 4049 -26
rect 4049 -288 4058 -26
rect 4006 -294 4058 -288
rect 4102 288 4154 294
rect 4102 26 4111 288
rect 4111 26 4145 288
rect 4145 26 4154 288
rect 4198 -288 4207 -26
rect 4207 -288 4241 -26
rect 4241 -288 4250 -26
rect 4198 -294 4250 -288
rect 4294 288 4346 294
rect 4294 26 4303 288
rect 4303 26 4337 288
rect 4337 26 4346 288
rect 4390 -288 4399 -26
rect 4399 -288 4433 -26
rect 4433 -288 4442 -26
rect 4390 -294 4442 -288
rect 4486 288 4538 294
rect 4486 26 4495 288
rect 4495 26 4529 288
rect 4529 26 4538 288
rect 4582 -288 4591 -26
rect 4591 -288 4625 -26
rect 4625 -288 4634 -26
rect 4582 -294 4634 -288
rect 4678 288 4730 294
rect 4678 26 4687 288
rect 4687 26 4721 288
rect 4721 26 4730 288
rect 4774 -288 4783 -26
rect 4783 -288 4817 -26
rect 4817 -288 4826 -26
rect 4774 -294 4826 -288
rect 4870 288 4922 294
rect 4870 26 4879 288
rect 4879 26 4913 288
rect 4913 26 4922 288
rect 4966 -288 4975 -26
rect 4975 -288 5009 -26
rect 5009 -288 5018 -26
rect 4966 -294 5018 -288
rect 5062 288 5114 294
rect 5062 26 5071 288
rect 5071 26 5105 288
rect 5105 26 5114 288
rect 5158 -288 5167 -26
rect 5167 -288 5201 -26
rect 5201 -288 5210 -26
rect 5158 -294 5210 -288
rect 5254 288 5306 294
rect 5254 26 5263 288
rect 5263 26 5297 288
rect 5297 26 5306 288
rect 5350 -288 5359 -26
rect 5359 -288 5393 -26
rect 5393 -288 5402 -26
rect 5350 -294 5402 -288
rect 5446 288 5498 294
rect 5446 26 5455 288
rect 5455 26 5489 288
rect 5489 26 5498 288
rect 5542 -288 5551 -26
rect 5551 -288 5585 -26
rect 5585 -288 5594 -26
rect 5542 -294 5594 -288
rect 5638 288 5690 294
rect 5638 26 5647 288
rect 5647 26 5681 288
rect 5681 26 5690 288
rect 5734 -288 5743 -26
rect 5743 -288 5777 -26
rect 5777 -288 5786 -26
rect 5734 -294 5786 -288
<< metal2 >>
rect -5690 294 5690 300
rect -5638 26 -5498 294
rect -5446 26 -5306 294
rect -5254 26 -5114 294
rect -5062 26 -4922 294
rect -4870 26 -4730 294
rect -4678 26 -4538 294
rect -4486 26 -4346 294
rect -4294 26 -4154 294
rect -4102 26 -3962 294
rect -3910 26 -3770 294
rect -3718 26 -3578 294
rect -3526 26 -3386 294
rect -3334 26 -3194 294
rect -3142 26 -3002 294
rect -2950 26 -2810 294
rect -2758 26 -2618 294
rect -2566 26 -2426 294
rect -2374 26 -2234 294
rect -2182 26 -2042 294
rect -1990 26 -1850 294
rect -1798 26 -1658 294
rect -1606 26 -1466 294
rect -1414 26 -1274 294
rect -1222 26 -1082 294
rect -1030 26 -890 294
rect -838 26 -698 294
rect -646 26 -506 294
rect -454 26 -314 294
rect -262 26 -122 294
rect -70 26 70 294
rect 122 26 262 294
rect 314 26 454 294
rect 506 26 646 294
rect 698 26 838 294
rect 890 26 1030 294
rect 1082 26 1222 294
rect 1274 26 1414 294
rect 1466 26 1606 294
rect 1658 26 1798 294
rect 1850 26 1990 294
rect 2042 26 2182 294
rect 2234 26 2374 294
rect 2426 26 2566 294
rect 2618 26 2758 294
rect 2810 26 2950 294
rect 3002 26 3142 294
rect 3194 26 3334 294
rect 3386 26 3526 294
rect 3578 26 3718 294
rect 3770 26 3910 294
rect 3962 26 4102 294
rect 4154 26 4294 294
rect 4346 26 4486 294
rect 4538 26 4678 294
rect 4730 26 4870 294
rect 4922 26 5062 294
rect 5114 26 5254 294
rect 5306 26 5446 294
rect 5498 26 5638 294
rect -5690 20 5690 26
rect -5786 -26 5786 -20
rect -5734 -294 -5594 -26
rect -5542 -294 -5402 -26
rect -5350 -294 -5210 -26
rect -5158 -294 -5018 -26
rect -4966 -294 -4826 -26
rect -4774 -294 -4634 -26
rect -4582 -294 -4442 -26
rect -4390 -294 -4250 -26
rect -4198 -294 -4058 -26
rect -4006 -294 -3866 -26
rect -3814 -294 -3674 -26
rect -3622 -294 -3482 -26
rect -3430 -294 -3290 -26
rect -3238 -294 -3098 -26
rect -3046 -294 -2906 -26
rect -2854 -294 -2714 -26
rect -2662 -294 -2522 -26
rect -2470 -294 -2330 -26
rect -2278 -294 -2138 -26
rect -2086 -294 -1946 -26
rect -1894 -294 -1754 -26
rect -1702 -294 -1562 -26
rect -1510 -294 -1370 -26
rect -1318 -294 -1178 -26
rect -1126 -294 -986 -26
rect -934 -294 -794 -26
rect -742 -294 -602 -26
rect -550 -294 -410 -26
rect -358 -294 -218 -26
rect -166 -294 -26 -26
rect 26 -294 166 -26
rect 218 -294 358 -26
rect 410 -294 550 -26
rect 602 -294 742 -26
rect 794 -294 934 -26
rect 986 -294 1126 -26
rect 1178 -294 1318 -26
rect 1370 -294 1510 -26
rect 1562 -294 1702 -26
rect 1754 -294 1894 -26
rect 1946 -294 2086 -26
rect 2138 -294 2278 -26
rect 2330 -294 2470 -26
rect 2522 -294 2662 -26
rect 2714 -294 2854 -26
rect 2906 -294 3046 -26
rect 3098 -294 3238 -26
rect 3290 -294 3430 -26
rect 3482 -294 3622 -26
rect 3674 -294 3814 -26
rect 3866 -294 4006 -26
rect 4058 -294 4198 -26
rect 4250 -294 4390 -26
rect 4442 -294 4582 -26
rect 4634 -294 4774 -26
rect 4826 -294 4966 -26
rect 5018 -294 5158 -26
rect 5210 -294 5350 -26
rect 5402 -294 5542 -26
rect 5594 -294 5734 -26
rect -5786 -300 5786 -294
<< properties >>
string FIXED_BBOX -5874 -466 5874 466
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 3 l 0.15 m 1 nf 120 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
