magic
tech sky130A
magscale 1 2
timestamp 1725098041
<< nwell >>
rect -6549 -597 6549 597
<< mvpmos >>
rect -6291 -300 -6191 300
rect -6133 -300 -6033 300
rect -5975 -300 -5875 300
rect -5817 -300 -5717 300
rect -5659 -300 -5559 300
rect -5501 -300 -5401 300
rect -5343 -300 -5243 300
rect -5185 -300 -5085 300
rect -5027 -300 -4927 300
rect -4869 -300 -4769 300
rect -4711 -300 -4611 300
rect -4553 -300 -4453 300
rect -4395 -300 -4295 300
rect -4237 -300 -4137 300
rect -4079 -300 -3979 300
rect -3921 -300 -3821 300
rect -3763 -300 -3663 300
rect -3605 -300 -3505 300
rect -3447 -300 -3347 300
rect -3289 -300 -3189 300
rect -3131 -300 -3031 300
rect -2973 -300 -2873 300
rect -2815 -300 -2715 300
rect -2657 -300 -2557 300
rect -2499 -300 -2399 300
rect -2341 -300 -2241 300
rect -2183 -300 -2083 300
rect -2025 -300 -1925 300
rect -1867 -300 -1767 300
rect -1709 -300 -1609 300
rect -1551 -300 -1451 300
rect -1393 -300 -1293 300
rect -1235 -300 -1135 300
rect -1077 -300 -977 300
rect -919 -300 -819 300
rect -761 -300 -661 300
rect -603 -300 -503 300
rect -445 -300 -345 300
rect -287 -300 -187 300
rect -129 -300 -29 300
rect 29 -300 129 300
rect 187 -300 287 300
rect 345 -300 445 300
rect 503 -300 603 300
rect 661 -300 761 300
rect 819 -300 919 300
rect 977 -300 1077 300
rect 1135 -300 1235 300
rect 1293 -300 1393 300
rect 1451 -300 1551 300
rect 1609 -300 1709 300
rect 1767 -300 1867 300
rect 1925 -300 2025 300
rect 2083 -300 2183 300
rect 2241 -300 2341 300
rect 2399 -300 2499 300
rect 2557 -300 2657 300
rect 2715 -300 2815 300
rect 2873 -300 2973 300
rect 3031 -300 3131 300
rect 3189 -300 3289 300
rect 3347 -300 3447 300
rect 3505 -300 3605 300
rect 3663 -300 3763 300
rect 3821 -300 3921 300
rect 3979 -300 4079 300
rect 4137 -300 4237 300
rect 4295 -300 4395 300
rect 4453 -300 4553 300
rect 4611 -300 4711 300
rect 4769 -300 4869 300
rect 4927 -300 5027 300
rect 5085 -300 5185 300
rect 5243 -300 5343 300
rect 5401 -300 5501 300
rect 5559 -300 5659 300
rect 5717 -300 5817 300
rect 5875 -300 5975 300
rect 6033 -300 6133 300
rect 6191 -300 6291 300
<< mvpdiff >>
rect -6349 288 -6291 300
rect -6349 -288 -6337 288
rect -6303 -288 -6291 288
rect -6349 -300 -6291 -288
rect -6191 288 -6133 300
rect -6191 -288 -6179 288
rect -6145 -288 -6133 288
rect -6191 -300 -6133 -288
rect -6033 288 -5975 300
rect -6033 -288 -6021 288
rect -5987 -288 -5975 288
rect -6033 -300 -5975 -288
rect -5875 288 -5817 300
rect -5875 -288 -5863 288
rect -5829 -288 -5817 288
rect -5875 -300 -5817 -288
rect -5717 288 -5659 300
rect -5717 -288 -5705 288
rect -5671 -288 -5659 288
rect -5717 -300 -5659 -288
rect -5559 288 -5501 300
rect -5559 -288 -5547 288
rect -5513 -288 -5501 288
rect -5559 -300 -5501 -288
rect -5401 288 -5343 300
rect -5401 -288 -5389 288
rect -5355 -288 -5343 288
rect -5401 -300 -5343 -288
rect -5243 288 -5185 300
rect -5243 -288 -5231 288
rect -5197 -288 -5185 288
rect -5243 -300 -5185 -288
rect -5085 288 -5027 300
rect -5085 -288 -5073 288
rect -5039 -288 -5027 288
rect -5085 -300 -5027 -288
rect -4927 288 -4869 300
rect -4927 -288 -4915 288
rect -4881 -288 -4869 288
rect -4927 -300 -4869 -288
rect -4769 288 -4711 300
rect -4769 -288 -4757 288
rect -4723 -288 -4711 288
rect -4769 -300 -4711 -288
rect -4611 288 -4553 300
rect -4611 -288 -4599 288
rect -4565 -288 -4553 288
rect -4611 -300 -4553 -288
rect -4453 288 -4395 300
rect -4453 -288 -4441 288
rect -4407 -288 -4395 288
rect -4453 -300 -4395 -288
rect -4295 288 -4237 300
rect -4295 -288 -4283 288
rect -4249 -288 -4237 288
rect -4295 -300 -4237 -288
rect -4137 288 -4079 300
rect -4137 -288 -4125 288
rect -4091 -288 -4079 288
rect -4137 -300 -4079 -288
rect -3979 288 -3921 300
rect -3979 -288 -3967 288
rect -3933 -288 -3921 288
rect -3979 -300 -3921 -288
rect -3821 288 -3763 300
rect -3821 -288 -3809 288
rect -3775 -288 -3763 288
rect -3821 -300 -3763 -288
rect -3663 288 -3605 300
rect -3663 -288 -3651 288
rect -3617 -288 -3605 288
rect -3663 -300 -3605 -288
rect -3505 288 -3447 300
rect -3505 -288 -3493 288
rect -3459 -288 -3447 288
rect -3505 -300 -3447 -288
rect -3347 288 -3289 300
rect -3347 -288 -3335 288
rect -3301 -288 -3289 288
rect -3347 -300 -3289 -288
rect -3189 288 -3131 300
rect -3189 -288 -3177 288
rect -3143 -288 -3131 288
rect -3189 -300 -3131 -288
rect -3031 288 -2973 300
rect -3031 -288 -3019 288
rect -2985 -288 -2973 288
rect -3031 -300 -2973 -288
rect -2873 288 -2815 300
rect -2873 -288 -2861 288
rect -2827 -288 -2815 288
rect -2873 -300 -2815 -288
rect -2715 288 -2657 300
rect -2715 -288 -2703 288
rect -2669 -288 -2657 288
rect -2715 -300 -2657 -288
rect -2557 288 -2499 300
rect -2557 -288 -2545 288
rect -2511 -288 -2499 288
rect -2557 -300 -2499 -288
rect -2399 288 -2341 300
rect -2399 -288 -2387 288
rect -2353 -288 -2341 288
rect -2399 -300 -2341 -288
rect -2241 288 -2183 300
rect -2241 -288 -2229 288
rect -2195 -288 -2183 288
rect -2241 -300 -2183 -288
rect -2083 288 -2025 300
rect -2083 -288 -2071 288
rect -2037 -288 -2025 288
rect -2083 -300 -2025 -288
rect -1925 288 -1867 300
rect -1925 -288 -1913 288
rect -1879 -288 -1867 288
rect -1925 -300 -1867 -288
rect -1767 288 -1709 300
rect -1767 -288 -1755 288
rect -1721 -288 -1709 288
rect -1767 -300 -1709 -288
rect -1609 288 -1551 300
rect -1609 -288 -1597 288
rect -1563 -288 -1551 288
rect -1609 -300 -1551 -288
rect -1451 288 -1393 300
rect -1451 -288 -1439 288
rect -1405 -288 -1393 288
rect -1451 -300 -1393 -288
rect -1293 288 -1235 300
rect -1293 -288 -1281 288
rect -1247 -288 -1235 288
rect -1293 -300 -1235 -288
rect -1135 288 -1077 300
rect -1135 -288 -1123 288
rect -1089 -288 -1077 288
rect -1135 -300 -1077 -288
rect -977 288 -919 300
rect -977 -288 -965 288
rect -931 -288 -919 288
rect -977 -300 -919 -288
rect -819 288 -761 300
rect -819 -288 -807 288
rect -773 -288 -761 288
rect -819 -300 -761 -288
rect -661 288 -603 300
rect -661 -288 -649 288
rect -615 -288 -603 288
rect -661 -300 -603 -288
rect -503 288 -445 300
rect -503 -288 -491 288
rect -457 -288 -445 288
rect -503 -300 -445 -288
rect -345 288 -287 300
rect -345 -288 -333 288
rect -299 -288 -287 288
rect -345 -300 -287 -288
rect -187 288 -129 300
rect -187 -288 -175 288
rect -141 -288 -129 288
rect -187 -300 -129 -288
rect -29 288 29 300
rect -29 -288 -17 288
rect 17 -288 29 288
rect -29 -300 29 -288
rect 129 288 187 300
rect 129 -288 141 288
rect 175 -288 187 288
rect 129 -300 187 -288
rect 287 288 345 300
rect 287 -288 299 288
rect 333 -288 345 288
rect 287 -300 345 -288
rect 445 288 503 300
rect 445 -288 457 288
rect 491 -288 503 288
rect 445 -300 503 -288
rect 603 288 661 300
rect 603 -288 615 288
rect 649 -288 661 288
rect 603 -300 661 -288
rect 761 288 819 300
rect 761 -288 773 288
rect 807 -288 819 288
rect 761 -300 819 -288
rect 919 288 977 300
rect 919 -288 931 288
rect 965 -288 977 288
rect 919 -300 977 -288
rect 1077 288 1135 300
rect 1077 -288 1089 288
rect 1123 -288 1135 288
rect 1077 -300 1135 -288
rect 1235 288 1293 300
rect 1235 -288 1247 288
rect 1281 -288 1293 288
rect 1235 -300 1293 -288
rect 1393 288 1451 300
rect 1393 -288 1405 288
rect 1439 -288 1451 288
rect 1393 -300 1451 -288
rect 1551 288 1609 300
rect 1551 -288 1563 288
rect 1597 -288 1609 288
rect 1551 -300 1609 -288
rect 1709 288 1767 300
rect 1709 -288 1721 288
rect 1755 -288 1767 288
rect 1709 -300 1767 -288
rect 1867 288 1925 300
rect 1867 -288 1879 288
rect 1913 -288 1925 288
rect 1867 -300 1925 -288
rect 2025 288 2083 300
rect 2025 -288 2037 288
rect 2071 -288 2083 288
rect 2025 -300 2083 -288
rect 2183 288 2241 300
rect 2183 -288 2195 288
rect 2229 -288 2241 288
rect 2183 -300 2241 -288
rect 2341 288 2399 300
rect 2341 -288 2353 288
rect 2387 -288 2399 288
rect 2341 -300 2399 -288
rect 2499 288 2557 300
rect 2499 -288 2511 288
rect 2545 -288 2557 288
rect 2499 -300 2557 -288
rect 2657 288 2715 300
rect 2657 -288 2669 288
rect 2703 -288 2715 288
rect 2657 -300 2715 -288
rect 2815 288 2873 300
rect 2815 -288 2827 288
rect 2861 -288 2873 288
rect 2815 -300 2873 -288
rect 2973 288 3031 300
rect 2973 -288 2985 288
rect 3019 -288 3031 288
rect 2973 -300 3031 -288
rect 3131 288 3189 300
rect 3131 -288 3143 288
rect 3177 -288 3189 288
rect 3131 -300 3189 -288
rect 3289 288 3347 300
rect 3289 -288 3301 288
rect 3335 -288 3347 288
rect 3289 -300 3347 -288
rect 3447 288 3505 300
rect 3447 -288 3459 288
rect 3493 -288 3505 288
rect 3447 -300 3505 -288
rect 3605 288 3663 300
rect 3605 -288 3617 288
rect 3651 -288 3663 288
rect 3605 -300 3663 -288
rect 3763 288 3821 300
rect 3763 -288 3775 288
rect 3809 -288 3821 288
rect 3763 -300 3821 -288
rect 3921 288 3979 300
rect 3921 -288 3933 288
rect 3967 -288 3979 288
rect 3921 -300 3979 -288
rect 4079 288 4137 300
rect 4079 -288 4091 288
rect 4125 -288 4137 288
rect 4079 -300 4137 -288
rect 4237 288 4295 300
rect 4237 -288 4249 288
rect 4283 -288 4295 288
rect 4237 -300 4295 -288
rect 4395 288 4453 300
rect 4395 -288 4407 288
rect 4441 -288 4453 288
rect 4395 -300 4453 -288
rect 4553 288 4611 300
rect 4553 -288 4565 288
rect 4599 -288 4611 288
rect 4553 -300 4611 -288
rect 4711 288 4769 300
rect 4711 -288 4723 288
rect 4757 -288 4769 288
rect 4711 -300 4769 -288
rect 4869 288 4927 300
rect 4869 -288 4881 288
rect 4915 -288 4927 288
rect 4869 -300 4927 -288
rect 5027 288 5085 300
rect 5027 -288 5039 288
rect 5073 -288 5085 288
rect 5027 -300 5085 -288
rect 5185 288 5243 300
rect 5185 -288 5197 288
rect 5231 -288 5243 288
rect 5185 -300 5243 -288
rect 5343 288 5401 300
rect 5343 -288 5355 288
rect 5389 -288 5401 288
rect 5343 -300 5401 -288
rect 5501 288 5559 300
rect 5501 -288 5513 288
rect 5547 -288 5559 288
rect 5501 -300 5559 -288
rect 5659 288 5717 300
rect 5659 -288 5671 288
rect 5705 -288 5717 288
rect 5659 -300 5717 -288
rect 5817 288 5875 300
rect 5817 -288 5829 288
rect 5863 -288 5875 288
rect 5817 -300 5875 -288
rect 5975 288 6033 300
rect 5975 -288 5987 288
rect 6021 -288 6033 288
rect 5975 -300 6033 -288
rect 6133 288 6191 300
rect 6133 -288 6145 288
rect 6179 -288 6191 288
rect 6133 -300 6191 -288
rect 6291 288 6349 300
rect 6291 -288 6303 288
rect 6337 -288 6349 288
rect 6291 -300 6349 -288
<< mvpdiffc >>
rect -6337 -288 -6303 288
rect -6179 -288 -6145 288
rect -6021 -288 -5987 288
rect -5863 -288 -5829 288
rect -5705 -288 -5671 288
rect -5547 -288 -5513 288
rect -5389 -288 -5355 288
rect -5231 -288 -5197 288
rect -5073 -288 -5039 288
rect -4915 -288 -4881 288
rect -4757 -288 -4723 288
rect -4599 -288 -4565 288
rect -4441 -288 -4407 288
rect -4283 -288 -4249 288
rect -4125 -288 -4091 288
rect -3967 -288 -3933 288
rect -3809 -288 -3775 288
rect -3651 -288 -3617 288
rect -3493 -288 -3459 288
rect -3335 -288 -3301 288
rect -3177 -288 -3143 288
rect -3019 -288 -2985 288
rect -2861 -288 -2827 288
rect -2703 -288 -2669 288
rect -2545 -288 -2511 288
rect -2387 -288 -2353 288
rect -2229 -288 -2195 288
rect -2071 -288 -2037 288
rect -1913 -288 -1879 288
rect -1755 -288 -1721 288
rect -1597 -288 -1563 288
rect -1439 -288 -1405 288
rect -1281 -288 -1247 288
rect -1123 -288 -1089 288
rect -965 -288 -931 288
rect -807 -288 -773 288
rect -649 -288 -615 288
rect -491 -288 -457 288
rect -333 -288 -299 288
rect -175 -288 -141 288
rect -17 -288 17 288
rect 141 -288 175 288
rect 299 -288 333 288
rect 457 -288 491 288
rect 615 -288 649 288
rect 773 -288 807 288
rect 931 -288 965 288
rect 1089 -288 1123 288
rect 1247 -288 1281 288
rect 1405 -288 1439 288
rect 1563 -288 1597 288
rect 1721 -288 1755 288
rect 1879 -288 1913 288
rect 2037 -288 2071 288
rect 2195 -288 2229 288
rect 2353 -288 2387 288
rect 2511 -288 2545 288
rect 2669 -288 2703 288
rect 2827 -288 2861 288
rect 2985 -288 3019 288
rect 3143 -288 3177 288
rect 3301 -288 3335 288
rect 3459 -288 3493 288
rect 3617 -288 3651 288
rect 3775 -288 3809 288
rect 3933 -288 3967 288
rect 4091 -288 4125 288
rect 4249 -288 4283 288
rect 4407 -288 4441 288
rect 4565 -288 4599 288
rect 4723 -288 4757 288
rect 4881 -288 4915 288
rect 5039 -288 5073 288
rect 5197 -288 5231 288
rect 5355 -288 5389 288
rect 5513 -288 5547 288
rect 5671 -288 5705 288
rect 5829 -288 5863 288
rect 5987 -288 6021 288
rect 6145 -288 6179 288
rect 6303 -288 6337 288
<< mvnsubdiff >>
rect -6483 519 6483 531
rect -6483 485 -6375 519
rect 6375 485 6483 519
rect -6483 473 6483 485
rect -6483 423 -6425 473
rect -6483 -423 -6471 423
rect -6437 -423 -6425 423
rect 6425 423 6483 473
rect -6483 -473 -6425 -423
rect 6425 -423 6437 423
rect 6471 -423 6483 423
rect 6425 -473 6483 -423
rect -6483 -485 6483 -473
rect -6483 -519 -6375 -485
rect 6375 -519 6483 -485
rect -6483 -531 6483 -519
<< mvnsubdiffcont >>
rect -6375 485 6375 519
rect -6471 -423 -6437 423
rect 6437 -423 6471 423
rect -6375 -519 6375 -485
<< poly >>
rect -6291 381 -6191 397
rect -6291 347 -6275 381
rect -6207 347 -6191 381
rect -6291 300 -6191 347
rect -6133 381 -6033 397
rect -6133 347 -6117 381
rect -6049 347 -6033 381
rect -6133 300 -6033 347
rect -5975 381 -5875 397
rect -5975 347 -5959 381
rect -5891 347 -5875 381
rect -5975 300 -5875 347
rect -5817 381 -5717 397
rect -5817 347 -5801 381
rect -5733 347 -5717 381
rect -5817 300 -5717 347
rect -5659 381 -5559 397
rect -5659 347 -5643 381
rect -5575 347 -5559 381
rect -5659 300 -5559 347
rect -5501 381 -5401 397
rect -5501 347 -5485 381
rect -5417 347 -5401 381
rect -5501 300 -5401 347
rect -5343 381 -5243 397
rect -5343 347 -5327 381
rect -5259 347 -5243 381
rect -5343 300 -5243 347
rect -5185 381 -5085 397
rect -5185 347 -5169 381
rect -5101 347 -5085 381
rect -5185 300 -5085 347
rect -5027 381 -4927 397
rect -5027 347 -5011 381
rect -4943 347 -4927 381
rect -5027 300 -4927 347
rect -4869 381 -4769 397
rect -4869 347 -4853 381
rect -4785 347 -4769 381
rect -4869 300 -4769 347
rect -4711 381 -4611 397
rect -4711 347 -4695 381
rect -4627 347 -4611 381
rect -4711 300 -4611 347
rect -4553 381 -4453 397
rect -4553 347 -4537 381
rect -4469 347 -4453 381
rect -4553 300 -4453 347
rect -4395 381 -4295 397
rect -4395 347 -4379 381
rect -4311 347 -4295 381
rect -4395 300 -4295 347
rect -4237 381 -4137 397
rect -4237 347 -4221 381
rect -4153 347 -4137 381
rect -4237 300 -4137 347
rect -4079 381 -3979 397
rect -4079 347 -4063 381
rect -3995 347 -3979 381
rect -4079 300 -3979 347
rect -3921 381 -3821 397
rect -3921 347 -3905 381
rect -3837 347 -3821 381
rect -3921 300 -3821 347
rect -3763 381 -3663 397
rect -3763 347 -3747 381
rect -3679 347 -3663 381
rect -3763 300 -3663 347
rect -3605 381 -3505 397
rect -3605 347 -3589 381
rect -3521 347 -3505 381
rect -3605 300 -3505 347
rect -3447 381 -3347 397
rect -3447 347 -3431 381
rect -3363 347 -3347 381
rect -3447 300 -3347 347
rect -3289 381 -3189 397
rect -3289 347 -3273 381
rect -3205 347 -3189 381
rect -3289 300 -3189 347
rect -3131 381 -3031 397
rect -3131 347 -3115 381
rect -3047 347 -3031 381
rect -3131 300 -3031 347
rect -2973 381 -2873 397
rect -2973 347 -2957 381
rect -2889 347 -2873 381
rect -2973 300 -2873 347
rect -2815 381 -2715 397
rect -2815 347 -2799 381
rect -2731 347 -2715 381
rect -2815 300 -2715 347
rect -2657 381 -2557 397
rect -2657 347 -2641 381
rect -2573 347 -2557 381
rect -2657 300 -2557 347
rect -2499 381 -2399 397
rect -2499 347 -2483 381
rect -2415 347 -2399 381
rect -2499 300 -2399 347
rect -2341 381 -2241 397
rect -2341 347 -2325 381
rect -2257 347 -2241 381
rect -2341 300 -2241 347
rect -2183 381 -2083 397
rect -2183 347 -2167 381
rect -2099 347 -2083 381
rect -2183 300 -2083 347
rect -2025 381 -1925 397
rect -2025 347 -2009 381
rect -1941 347 -1925 381
rect -2025 300 -1925 347
rect -1867 381 -1767 397
rect -1867 347 -1851 381
rect -1783 347 -1767 381
rect -1867 300 -1767 347
rect -1709 381 -1609 397
rect -1709 347 -1693 381
rect -1625 347 -1609 381
rect -1709 300 -1609 347
rect -1551 381 -1451 397
rect -1551 347 -1535 381
rect -1467 347 -1451 381
rect -1551 300 -1451 347
rect -1393 381 -1293 397
rect -1393 347 -1377 381
rect -1309 347 -1293 381
rect -1393 300 -1293 347
rect -1235 381 -1135 397
rect -1235 347 -1219 381
rect -1151 347 -1135 381
rect -1235 300 -1135 347
rect -1077 381 -977 397
rect -1077 347 -1061 381
rect -993 347 -977 381
rect -1077 300 -977 347
rect -919 381 -819 397
rect -919 347 -903 381
rect -835 347 -819 381
rect -919 300 -819 347
rect -761 381 -661 397
rect -761 347 -745 381
rect -677 347 -661 381
rect -761 300 -661 347
rect -603 381 -503 397
rect -603 347 -587 381
rect -519 347 -503 381
rect -603 300 -503 347
rect -445 381 -345 397
rect -445 347 -429 381
rect -361 347 -345 381
rect -445 300 -345 347
rect -287 381 -187 397
rect -287 347 -271 381
rect -203 347 -187 381
rect -287 300 -187 347
rect -129 381 -29 397
rect -129 347 -113 381
rect -45 347 -29 381
rect -129 300 -29 347
rect 29 381 129 397
rect 29 347 45 381
rect 113 347 129 381
rect 29 300 129 347
rect 187 381 287 397
rect 187 347 203 381
rect 271 347 287 381
rect 187 300 287 347
rect 345 381 445 397
rect 345 347 361 381
rect 429 347 445 381
rect 345 300 445 347
rect 503 381 603 397
rect 503 347 519 381
rect 587 347 603 381
rect 503 300 603 347
rect 661 381 761 397
rect 661 347 677 381
rect 745 347 761 381
rect 661 300 761 347
rect 819 381 919 397
rect 819 347 835 381
rect 903 347 919 381
rect 819 300 919 347
rect 977 381 1077 397
rect 977 347 993 381
rect 1061 347 1077 381
rect 977 300 1077 347
rect 1135 381 1235 397
rect 1135 347 1151 381
rect 1219 347 1235 381
rect 1135 300 1235 347
rect 1293 381 1393 397
rect 1293 347 1309 381
rect 1377 347 1393 381
rect 1293 300 1393 347
rect 1451 381 1551 397
rect 1451 347 1467 381
rect 1535 347 1551 381
rect 1451 300 1551 347
rect 1609 381 1709 397
rect 1609 347 1625 381
rect 1693 347 1709 381
rect 1609 300 1709 347
rect 1767 381 1867 397
rect 1767 347 1783 381
rect 1851 347 1867 381
rect 1767 300 1867 347
rect 1925 381 2025 397
rect 1925 347 1941 381
rect 2009 347 2025 381
rect 1925 300 2025 347
rect 2083 381 2183 397
rect 2083 347 2099 381
rect 2167 347 2183 381
rect 2083 300 2183 347
rect 2241 381 2341 397
rect 2241 347 2257 381
rect 2325 347 2341 381
rect 2241 300 2341 347
rect 2399 381 2499 397
rect 2399 347 2415 381
rect 2483 347 2499 381
rect 2399 300 2499 347
rect 2557 381 2657 397
rect 2557 347 2573 381
rect 2641 347 2657 381
rect 2557 300 2657 347
rect 2715 381 2815 397
rect 2715 347 2731 381
rect 2799 347 2815 381
rect 2715 300 2815 347
rect 2873 381 2973 397
rect 2873 347 2889 381
rect 2957 347 2973 381
rect 2873 300 2973 347
rect 3031 381 3131 397
rect 3031 347 3047 381
rect 3115 347 3131 381
rect 3031 300 3131 347
rect 3189 381 3289 397
rect 3189 347 3205 381
rect 3273 347 3289 381
rect 3189 300 3289 347
rect 3347 381 3447 397
rect 3347 347 3363 381
rect 3431 347 3447 381
rect 3347 300 3447 347
rect 3505 381 3605 397
rect 3505 347 3521 381
rect 3589 347 3605 381
rect 3505 300 3605 347
rect 3663 381 3763 397
rect 3663 347 3679 381
rect 3747 347 3763 381
rect 3663 300 3763 347
rect 3821 381 3921 397
rect 3821 347 3837 381
rect 3905 347 3921 381
rect 3821 300 3921 347
rect 3979 381 4079 397
rect 3979 347 3995 381
rect 4063 347 4079 381
rect 3979 300 4079 347
rect 4137 381 4237 397
rect 4137 347 4153 381
rect 4221 347 4237 381
rect 4137 300 4237 347
rect 4295 381 4395 397
rect 4295 347 4311 381
rect 4379 347 4395 381
rect 4295 300 4395 347
rect 4453 381 4553 397
rect 4453 347 4469 381
rect 4537 347 4553 381
rect 4453 300 4553 347
rect 4611 381 4711 397
rect 4611 347 4627 381
rect 4695 347 4711 381
rect 4611 300 4711 347
rect 4769 381 4869 397
rect 4769 347 4785 381
rect 4853 347 4869 381
rect 4769 300 4869 347
rect 4927 381 5027 397
rect 4927 347 4943 381
rect 5011 347 5027 381
rect 4927 300 5027 347
rect 5085 381 5185 397
rect 5085 347 5101 381
rect 5169 347 5185 381
rect 5085 300 5185 347
rect 5243 381 5343 397
rect 5243 347 5259 381
rect 5327 347 5343 381
rect 5243 300 5343 347
rect 5401 381 5501 397
rect 5401 347 5417 381
rect 5485 347 5501 381
rect 5401 300 5501 347
rect 5559 381 5659 397
rect 5559 347 5575 381
rect 5643 347 5659 381
rect 5559 300 5659 347
rect 5717 381 5817 397
rect 5717 347 5733 381
rect 5801 347 5817 381
rect 5717 300 5817 347
rect 5875 381 5975 397
rect 5875 347 5891 381
rect 5959 347 5975 381
rect 5875 300 5975 347
rect 6033 381 6133 397
rect 6033 347 6049 381
rect 6117 347 6133 381
rect 6033 300 6133 347
rect 6191 381 6291 397
rect 6191 347 6207 381
rect 6275 347 6291 381
rect 6191 300 6291 347
rect -6291 -347 -6191 -300
rect -6291 -381 -6275 -347
rect -6207 -381 -6191 -347
rect -6291 -397 -6191 -381
rect -6133 -347 -6033 -300
rect -6133 -381 -6117 -347
rect -6049 -381 -6033 -347
rect -6133 -397 -6033 -381
rect -5975 -347 -5875 -300
rect -5975 -381 -5959 -347
rect -5891 -381 -5875 -347
rect -5975 -397 -5875 -381
rect -5817 -347 -5717 -300
rect -5817 -381 -5801 -347
rect -5733 -381 -5717 -347
rect -5817 -397 -5717 -381
rect -5659 -347 -5559 -300
rect -5659 -381 -5643 -347
rect -5575 -381 -5559 -347
rect -5659 -397 -5559 -381
rect -5501 -347 -5401 -300
rect -5501 -381 -5485 -347
rect -5417 -381 -5401 -347
rect -5501 -397 -5401 -381
rect -5343 -347 -5243 -300
rect -5343 -381 -5327 -347
rect -5259 -381 -5243 -347
rect -5343 -397 -5243 -381
rect -5185 -347 -5085 -300
rect -5185 -381 -5169 -347
rect -5101 -381 -5085 -347
rect -5185 -397 -5085 -381
rect -5027 -347 -4927 -300
rect -5027 -381 -5011 -347
rect -4943 -381 -4927 -347
rect -5027 -397 -4927 -381
rect -4869 -347 -4769 -300
rect -4869 -381 -4853 -347
rect -4785 -381 -4769 -347
rect -4869 -397 -4769 -381
rect -4711 -347 -4611 -300
rect -4711 -381 -4695 -347
rect -4627 -381 -4611 -347
rect -4711 -397 -4611 -381
rect -4553 -347 -4453 -300
rect -4553 -381 -4537 -347
rect -4469 -381 -4453 -347
rect -4553 -397 -4453 -381
rect -4395 -347 -4295 -300
rect -4395 -381 -4379 -347
rect -4311 -381 -4295 -347
rect -4395 -397 -4295 -381
rect -4237 -347 -4137 -300
rect -4237 -381 -4221 -347
rect -4153 -381 -4137 -347
rect -4237 -397 -4137 -381
rect -4079 -347 -3979 -300
rect -4079 -381 -4063 -347
rect -3995 -381 -3979 -347
rect -4079 -397 -3979 -381
rect -3921 -347 -3821 -300
rect -3921 -381 -3905 -347
rect -3837 -381 -3821 -347
rect -3921 -397 -3821 -381
rect -3763 -347 -3663 -300
rect -3763 -381 -3747 -347
rect -3679 -381 -3663 -347
rect -3763 -397 -3663 -381
rect -3605 -347 -3505 -300
rect -3605 -381 -3589 -347
rect -3521 -381 -3505 -347
rect -3605 -397 -3505 -381
rect -3447 -347 -3347 -300
rect -3447 -381 -3431 -347
rect -3363 -381 -3347 -347
rect -3447 -397 -3347 -381
rect -3289 -347 -3189 -300
rect -3289 -381 -3273 -347
rect -3205 -381 -3189 -347
rect -3289 -397 -3189 -381
rect -3131 -347 -3031 -300
rect -3131 -381 -3115 -347
rect -3047 -381 -3031 -347
rect -3131 -397 -3031 -381
rect -2973 -347 -2873 -300
rect -2973 -381 -2957 -347
rect -2889 -381 -2873 -347
rect -2973 -397 -2873 -381
rect -2815 -347 -2715 -300
rect -2815 -381 -2799 -347
rect -2731 -381 -2715 -347
rect -2815 -397 -2715 -381
rect -2657 -347 -2557 -300
rect -2657 -381 -2641 -347
rect -2573 -381 -2557 -347
rect -2657 -397 -2557 -381
rect -2499 -347 -2399 -300
rect -2499 -381 -2483 -347
rect -2415 -381 -2399 -347
rect -2499 -397 -2399 -381
rect -2341 -347 -2241 -300
rect -2341 -381 -2325 -347
rect -2257 -381 -2241 -347
rect -2341 -397 -2241 -381
rect -2183 -347 -2083 -300
rect -2183 -381 -2167 -347
rect -2099 -381 -2083 -347
rect -2183 -397 -2083 -381
rect -2025 -347 -1925 -300
rect -2025 -381 -2009 -347
rect -1941 -381 -1925 -347
rect -2025 -397 -1925 -381
rect -1867 -347 -1767 -300
rect -1867 -381 -1851 -347
rect -1783 -381 -1767 -347
rect -1867 -397 -1767 -381
rect -1709 -347 -1609 -300
rect -1709 -381 -1693 -347
rect -1625 -381 -1609 -347
rect -1709 -397 -1609 -381
rect -1551 -347 -1451 -300
rect -1551 -381 -1535 -347
rect -1467 -381 -1451 -347
rect -1551 -397 -1451 -381
rect -1393 -347 -1293 -300
rect -1393 -381 -1377 -347
rect -1309 -381 -1293 -347
rect -1393 -397 -1293 -381
rect -1235 -347 -1135 -300
rect -1235 -381 -1219 -347
rect -1151 -381 -1135 -347
rect -1235 -397 -1135 -381
rect -1077 -347 -977 -300
rect -1077 -381 -1061 -347
rect -993 -381 -977 -347
rect -1077 -397 -977 -381
rect -919 -347 -819 -300
rect -919 -381 -903 -347
rect -835 -381 -819 -347
rect -919 -397 -819 -381
rect -761 -347 -661 -300
rect -761 -381 -745 -347
rect -677 -381 -661 -347
rect -761 -397 -661 -381
rect -603 -347 -503 -300
rect -603 -381 -587 -347
rect -519 -381 -503 -347
rect -603 -397 -503 -381
rect -445 -347 -345 -300
rect -445 -381 -429 -347
rect -361 -381 -345 -347
rect -445 -397 -345 -381
rect -287 -347 -187 -300
rect -287 -381 -271 -347
rect -203 -381 -187 -347
rect -287 -397 -187 -381
rect -129 -347 -29 -300
rect -129 -381 -113 -347
rect -45 -381 -29 -347
rect -129 -397 -29 -381
rect 29 -347 129 -300
rect 29 -381 45 -347
rect 113 -381 129 -347
rect 29 -397 129 -381
rect 187 -347 287 -300
rect 187 -381 203 -347
rect 271 -381 287 -347
rect 187 -397 287 -381
rect 345 -347 445 -300
rect 345 -381 361 -347
rect 429 -381 445 -347
rect 345 -397 445 -381
rect 503 -347 603 -300
rect 503 -381 519 -347
rect 587 -381 603 -347
rect 503 -397 603 -381
rect 661 -347 761 -300
rect 661 -381 677 -347
rect 745 -381 761 -347
rect 661 -397 761 -381
rect 819 -347 919 -300
rect 819 -381 835 -347
rect 903 -381 919 -347
rect 819 -397 919 -381
rect 977 -347 1077 -300
rect 977 -381 993 -347
rect 1061 -381 1077 -347
rect 977 -397 1077 -381
rect 1135 -347 1235 -300
rect 1135 -381 1151 -347
rect 1219 -381 1235 -347
rect 1135 -397 1235 -381
rect 1293 -347 1393 -300
rect 1293 -381 1309 -347
rect 1377 -381 1393 -347
rect 1293 -397 1393 -381
rect 1451 -347 1551 -300
rect 1451 -381 1467 -347
rect 1535 -381 1551 -347
rect 1451 -397 1551 -381
rect 1609 -347 1709 -300
rect 1609 -381 1625 -347
rect 1693 -381 1709 -347
rect 1609 -397 1709 -381
rect 1767 -347 1867 -300
rect 1767 -381 1783 -347
rect 1851 -381 1867 -347
rect 1767 -397 1867 -381
rect 1925 -347 2025 -300
rect 1925 -381 1941 -347
rect 2009 -381 2025 -347
rect 1925 -397 2025 -381
rect 2083 -347 2183 -300
rect 2083 -381 2099 -347
rect 2167 -381 2183 -347
rect 2083 -397 2183 -381
rect 2241 -347 2341 -300
rect 2241 -381 2257 -347
rect 2325 -381 2341 -347
rect 2241 -397 2341 -381
rect 2399 -347 2499 -300
rect 2399 -381 2415 -347
rect 2483 -381 2499 -347
rect 2399 -397 2499 -381
rect 2557 -347 2657 -300
rect 2557 -381 2573 -347
rect 2641 -381 2657 -347
rect 2557 -397 2657 -381
rect 2715 -347 2815 -300
rect 2715 -381 2731 -347
rect 2799 -381 2815 -347
rect 2715 -397 2815 -381
rect 2873 -347 2973 -300
rect 2873 -381 2889 -347
rect 2957 -381 2973 -347
rect 2873 -397 2973 -381
rect 3031 -347 3131 -300
rect 3031 -381 3047 -347
rect 3115 -381 3131 -347
rect 3031 -397 3131 -381
rect 3189 -347 3289 -300
rect 3189 -381 3205 -347
rect 3273 -381 3289 -347
rect 3189 -397 3289 -381
rect 3347 -347 3447 -300
rect 3347 -381 3363 -347
rect 3431 -381 3447 -347
rect 3347 -397 3447 -381
rect 3505 -347 3605 -300
rect 3505 -381 3521 -347
rect 3589 -381 3605 -347
rect 3505 -397 3605 -381
rect 3663 -347 3763 -300
rect 3663 -381 3679 -347
rect 3747 -381 3763 -347
rect 3663 -397 3763 -381
rect 3821 -347 3921 -300
rect 3821 -381 3837 -347
rect 3905 -381 3921 -347
rect 3821 -397 3921 -381
rect 3979 -347 4079 -300
rect 3979 -381 3995 -347
rect 4063 -381 4079 -347
rect 3979 -397 4079 -381
rect 4137 -347 4237 -300
rect 4137 -381 4153 -347
rect 4221 -381 4237 -347
rect 4137 -397 4237 -381
rect 4295 -347 4395 -300
rect 4295 -381 4311 -347
rect 4379 -381 4395 -347
rect 4295 -397 4395 -381
rect 4453 -347 4553 -300
rect 4453 -381 4469 -347
rect 4537 -381 4553 -347
rect 4453 -397 4553 -381
rect 4611 -347 4711 -300
rect 4611 -381 4627 -347
rect 4695 -381 4711 -347
rect 4611 -397 4711 -381
rect 4769 -347 4869 -300
rect 4769 -381 4785 -347
rect 4853 -381 4869 -347
rect 4769 -397 4869 -381
rect 4927 -347 5027 -300
rect 4927 -381 4943 -347
rect 5011 -381 5027 -347
rect 4927 -397 5027 -381
rect 5085 -347 5185 -300
rect 5085 -381 5101 -347
rect 5169 -381 5185 -347
rect 5085 -397 5185 -381
rect 5243 -347 5343 -300
rect 5243 -381 5259 -347
rect 5327 -381 5343 -347
rect 5243 -397 5343 -381
rect 5401 -347 5501 -300
rect 5401 -381 5417 -347
rect 5485 -381 5501 -347
rect 5401 -397 5501 -381
rect 5559 -347 5659 -300
rect 5559 -381 5575 -347
rect 5643 -381 5659 -347
rect 5559 -397 5659 -381
rect 5717 -347 5817 -300
rect 5717 -381 5733 -347
rect 5801 -381 5817 -347
rect 5717 -397 5817 -381
rect 5875 -347 5975 -300
rect 5875 -381 5891 -347
rect 5959 -381 5975 -347
rect 5875 -397 5975 -381
rect 6033 -347 6133 -300
rect 6033 -381 6049 -347
rect 6117 -381 6133 -347
rect 6033 -397 6133 -381
rect 6191 -347 6291 -300
rect 6191 -381 6207 -347
rect 6275 -381 6291 -347
rect 6191 -397 6291 -381
<< polycont >>
rect -6275 347 -6207 381
rect -6117 347 -6049 381
rect -5959 347 -5891 381
rect -5801 347 -5733 381
rect -5643 347 -5575 381
rect -5485 347 -5417 381
rect -5327 347 -5259 381
rect -5169 347 -5101 381
rect -5011 347 -4943 381
rect -4853 347 -4785 381
rect -4695 347 -4627 381
rect -4537 347 -4469 381
rect -4379 347 -4311 381
rect -4221 347 -4153 381
rect -4063 347 -3995 381
rect -3905 347 -3837 381
rect -3747 347 -3679 381
rect -3589 347 -3521 381
rect -3431 347 -3363 381
rect -3273 347 -3205 381
rect -3115 347 -3047 381
rect -2957 347 -2889 381
rect -2799 347 -2731 381
rect -2641 347 -2573 381
rect -2483 347 -2415 381
rect -2325 347 -2257 381
rect -2167 347 -2099 381
rect -2009 347 -1941 381
rect -1851 347 -1783 381
rect -1693 347 -1625 381
rect -1535 347 -1467 381
rect -1377 347 -1309 381
rect -1219 347 -1151 381
rect -1061 347 -993 381
rect -903 347 -835 381
rect -745 347 -677 381
rect -587 347 -519 381
rect -429 347 -361 381
rect -271 347 -203 381
rect -113 347 -45 381
rect 45 347 113 381
rect 203 347 271 381
rect 361 347 429 381
rect 519 347 587 381
rect 677 347 745 381
rect 835 347 903 381
rect 993 347 1061 381
rect 1151 347 1219 381
rect 1309 347 1377 381
rect 1467 347 1535 381
rect 1625 347 1693 381
rect 1783 347 1851 381
rect 1941 347 2009 381
rect 2099 347 2167 381
rect 2257 347 2325 381
rect 2415 347 2483 381
rect 2573 347 2641 381
rect 2731 347 2799 381
rect 2889 347 2957 381
rect 3047 347 3115 381
rect 3205 347 3273 381
rect 3363 347 3431 381
rect 3521 347 3589 381
rect 3679 347 3747 381
rect 3837 347 3905 381
rect 3995 347 4063 381
rect 4153 347 4221 381
rect 4311 347 4379 381
rect 4469 347 4537 381
rect 4627 347 4695 381
rect 4785 347 4853 381
rect 4943 347 5011 381
rect 5101 347 5169 381
rect 5259 347 5327 381
rect 5417 347 5485 381
rect 5575 347 5643 381
rect 5733 347 5801 381
rect 5891 347 5959 381
rect 6049 347 6117 381
rect 6207 347 6275 381
rect -6275 -381 -6207 -347
rect -6117 -381 -6049 -347
rect -5959 -381 -5891 -347
rect -5801 -381 -5733 -347
rect -5643 -381 -5575 -347
rect -5485 -381 -5417 -347
rect -5327 -381 -5259 -347
rect -5169 -381 -5101 -347
rect -5011 -381 -4943 -347
rect -4853 -381 -4785 -347
rect -4695 -381 -4627 -347
rect -4537 -381 -4469 -347
rect -4379 -381 -4311 -347
rect -4221 -381 -4153 -347
rect -4063 -381 -3995 -347
rect -3905 -381 -3837 -347
rect -3747 -381 -3679 -347
rect -3589 -381 -3521 -347
rect -3431 -381 -3363 -347
rect -3273 -381 -3205 -347
rect -3115 -381 -3047 -347
rect -2957 -381 -2889 -347
rect -2799 -381 -2731 -347
rect -2641 -381 -2573 -347
rect -2483 -381 -2415 -347
rect -2325 -381 -2257 -347
rect -2167 -381 -2099 -347
rect -2009 -381 -1941 -347
rect -1851 -381 -1783 -347
rect -1693 -381 -1625 -347
rect -1535 -381 -1467 -347
rect -1377 -381 -1309 -347
rect -1219 -381 -1151 -347
rect -1061 -381 -993 -347
rect -903 -381 -835 -347
rect -745 -381 -677 -347
rect -587 -381 -519 -347
rect -429 -381 -361 -347
rect -271 -381 -203 -347
rect -113 -381 -45 -347
rect 45 -381 113 -347
rect 203 -381 271 -347
rect 361 -381 429 -347
rect 519 -381 587 -347
rect 677 -381 745 -347
rect 835 -381 903 -347
rect 993 -381 1061 -347
rect 1151 -381 1219 -347
rect 1309 -381 1377 -347
rect 1467 -381 1535 -347
rect 1625 -381 1693 -347
rect 1783 -381 1851 -347
rect 1941 -381 2009 -347
rect 2099 -381 2167 -347
rect 2257 -381 2325 -347
rect 2415 -381 2483 -347
rect 2573 -381 2641 -347
rect 2731 -381 2799 -347
rect 2889 -381 2957 -347
rect 3047 -381 3115 -347
rect 3205 -381 3273 -347
rect 3363 -381 3431 -347
rect 3521 -381 3589 -347
rect 3679 -381 3747 -347
rect 3837 -381 3905 -347
rect 3995 -381 4063 -347
rect 4153 -381 4221 -347
rect 4311 -381 4379 -347
rect 4469 -381 4537 -347
rect 4627 -381 4695 -347
rect 4785 -381 4853 -347
rect 4943 -381 5011 -347
rect 5101 -381 5169 -347
rect 5259 -381 5327 -347
rect 5417 -381 5485 -347
rect 5575 -381 5643 -347
rect 5733 -381 5801 -347
rect 5891 -381 5959 -347
rect 6049 -381 6117 -347
rect 6207 -381 6275 -347
<< locali >>
rect 6375 485 6471 519
rect -6471 423 -6437 485
rect 6437 423 6471 485
rect -6291 347 -6275 381
rect -6207 347 -6117 381
rect -6049 347 -5959 381
rect -5891 347 -5801 381
rect -5733 347 -5643 381
rect -5575 347 -5485 381
rect -5417 347 -5327 381
rect -5259 347 -5169 381
rect -5101 347 -5011 381
rect -4943 347 -4853 381
rect -4785 347 -4695 381
rect -4627 347 -4537 381
rect -4469 347 -4379 381
rect -4311 347 -4221 381
rect -4153 347 -4063 381
rect -3995 347 -3905 381
rect -3837 347 -3747 381
rect -3679 347 -3589 381
rect -3521 347 -3431 381
rect -3363 347 -3273 381
rect -3205 347 -3115 381
rect -3047 347 -2957 381
rect -2889 347 -2799 381
rect -2731 347 -2641 381
rect -2573 347 -2483 381
rect -2415 347 -2325 381
rect -2257 347 -2167 381
rect -2099 347 -2009 381
rect -1941 347 -1851 381
rect -1783 347 -1693 381
rect -1625 347 -1535 381
rect -1467 347 -1377 381
rect -1309 347 -1219 381
rect -1151 347 -1061 381
rect -993 347 -903 381
rect -835 347 -745 381
rect -677 347 -587 381
rect -519 347 -429 381
rect -361 347 -271 381
rect -203 347 -113 381
rect -45 347 45 381
rect 113 347 203 381
rect 271 347 361 381
rect 429 347 519 381
rect 587 347 677 381
rect 745 347 835 381
rect 903 347 993 381
rect 1061 347 1151 381
rect 1219 347 1309 381
rect 1377 347 1467 381
rect 1535 347 1625 381
rect 1693 347 1783 381
rect 1851 347 1941 381
rect 2009 347 2099 381
rect 2167 347 2257 381
rect 2325 347 2415 381
rect 2483 347 2573 381
rect 2641 347 2731 381
rect 2799 347 2889 381
rect 2957 347 3047 381
rect 3115 347 3205 381
rect 3273 347 3363 381
rect 3431 347 3521 381
rect 3589 347 3679 381
rect 3747 347 3837 381
rect 3905 347 3995 381
rect 4063 347 4153 381
rect 4221 347 4311 381
rect 4379 347 4469 381
rect 4537 347 4627 381
rect 4695 347 4785 381
rect 4853 347 4943 381
rect 5011 347 5101 381
rect 5169 347 5259 381
rect 5327 347 5417 381
rect 5485 347 5575 381
rect 5643 347 5733 381
rect 5801 347 5891 381
rect 5959 347 6049 381
rect 6117 347 6207 381
rect 6275 347 6291 381
rect -6337 288 -6303 304
rect -6337 -304 -6303 -288
rect -6179 288 -6145 304
rect -6179 -304 -6145 -288
rect -6021 288 -5987 304
rect -6021 -304 -5987 -288
rect -5863 288 -5829 304
rect -5863 -304 -5829 -288
rect -5705 288 -5671 304
rect -5705 -304 -5671 -288
rect -5547 288 -5513 304
rect -5547 -304 -5513 -288
rect -5389 288 -5355 304
rect -5389 -304 -5355 -288
rect -5231 288 -5197 304
rect -5231 -304 -5197 -288
rect -5073 288 -5039 304
rect -5073 -304 -5039 -288
rect -4915 288 -4881 304
rect -4915 -304 -4881 -288
rect -4757 288 -4723 304
rect -4757 -304 -4723 -288
rect -4599 288 -4565 304
rect -4599 -304 -4565 -288
rect -4441 288 -4407 304
rect -4441 -304 -4407 -288
rect -4283 288 -4249 304
rect -4283 -304 -4249 -288
rect -4125 288 -4091 304
rect -4125 -304 -4091 -288
rect -3967 288 -3933 304
rect -3967 -304 -3933 -288
rect -3809 288 -3775 304
rect -3809 -304 -3775 -288
rect -3651 288 -3617 304
rect -3651 -304 -3617 -288
rect -3493 288 -3459 304
rect -3493 -304 -3459 -288
rect -3335 288 -3301 304
rect -3335 -304 -3301 -288
rect -3177 288 -3143 304
rect -3177 -304 -3143 -288
rect -3019 288 -2985 304
rect -3019 -304 -2985 -288
rect -2861 288 -2827 304
rect -2861 -304 -2827 -288
rect -2703 288 -2669 304
rect -2703 -304 -2669 -288
rect -2545 288 -2511 304
rect -2545 -304 -2511 -288
rect -2387 288 -2353 304
rect -2387 -304 -2353 -288
rect -2229 288 -2195 304
rect -2229 -304 -2195 -288
rect -2071 288 -2037 304
rect -2071 -304 -2037 -288
rect -1913 288 -1879 304
rect -1913 -304 -1879 -288
rect -1755 288 -1721 304
rect -1755 -304 -1721 -288
rect -1597 288 -1563 304
rect -1597 -304 -1563 -288
rect -1439 288 -1405 304
rect -1439 -304 -1405 -288
rect -1281 288 -1247 304
rect -1281 -304 -1247 -288
rect -1123 288 -1089 304
rect -1123 -304 -1089 -288
rect -965 288 -931 304
rect -965 -304 -931 -288
rect -807 288 -773 304
rect -807 -304 -773 -288
rect -649 288 -615 304
rect -649 -304 -615 -288
rect -491 288 -457 304
rect -491 -304 -457 -288
rect -333 288 -299 304
rect -333 -304 -299 -288
rect -175 288 -141 304
rect -175 -304 -141 -288
rect -17 288 17 304
rect -17 -304 17 -288
rect 141 288 175 304
rect 141 -304 175 -288
rect 299 288 333 304
rect 299 -304 333 -288
rect 457 288 491 304
rect 457 -304 491 -288
rect 615 288 649 304
rect 615 -304 649 -288
rect 773 288 807 304
rect 773 -304 807 -288
rect 931 288 965 304
rect 931 -304 965 -288
rect 1089 288 1123 304
rect 1089 -304 1123 -288
rect 1247 288 1281 304
rect 1247 -304 1281 -288
rect 1405 288 1439 304
rect 1405 -304 1439 -288
rect 1563 288 1597 304
rect 1563 -304 1597 -288
rect 1721 288 1755 304
rect 1721 -304 1755 -288
rect 1879 288 1913 304
rect 1879 -304 1913 -288
rect 2037 288 2071 304
rect 2037 -304 2071 -288
rect 2195 288 2229 304
rect 2195 -304 2229 -288
rect 2353 288 2387 304
rect 2353 -304 2387 -288
rect 2511 288 2545 304
rect 2511 -304 2545 -288
rect 2669 288 2703 304
rect 2669 -304 2703 -288
rect 2827 288 2861 304
rect 2827 -304 2861 -288
rect 2985 288 3019 304
rect 2985 -304 3019 -288
rect 3143 288 3177 304
rect 3143 -304 3177 -288
rect 3301 288 3335 304
rect 3301 -304 3335 -288
rect 3459 288 3493 304
rect 3459 -304 3493 -288
rect 3617 288 3651 304
rect 3617 -304 3651 -288
rect 3775 288 3809 304
rect 3775 -304 3809 -288
rect 3933 288 3967 304
rect 3933 -304 3967 -288
rect 4091 288 4125 304
rect 4091 -304 4125 -288
rect 4249 288 4283 304
rect 4249 -304 4283 -288
rect 4407 288 4441 304
rect 4407 -304 4441 -288
rect 4565 288 4599 304
rect 4565 -304 4599 -288
rect 4723 288 4757 304
rect 4723 -304 4757 -288
rect 4881 288 4915 304
rect 4881 -304 4915 -288
rect 5039 288 5073 304
rect 5039 -304 5073 -288
rect 5197 288 5231 304
rect 5197 -304 5231 -288
rect 5355 288 5389 304
rect 5355 -304 5389 -288
rect 5513 288 5547 304
rect 5513 -304 5547 -288
rect 5671 288 5705 304
rect 5671 -304 5705 -288
rect 5829 288 5863 304
rect 5829 -304 5863 -288
rect 5987 288 6021 304
rect 5987 -304 6021 -288
rect 6145 288 6179 304
rect 6145 -304 6179 -288
rect 6303 288 6337 304
rect 6303 -304 6337 -288
rect -6291 -381 -6275 -347
rect -6207 -381 -6117 -347
rect -6049 -381 -5959 -347
rect -5891 -381 -5801 -347
rect -5733 -381 -5643 -347
rect -5575 -381 -5485 -347
rect -5417 -381 -5327 -347
rect -5259 -381 -5169 -347
rect -5101 -381 -5011 -347
rect -4943 -381 -4853 -347
rect -4785 -381 -4695 -347
rect -4627 -381 -4537 -347
rect -4469 -381 -4379 -347
rect -4311 -381 -4221 -347
rect -4153 -381 -4063 -347
rect -3995 -381 -3905 -347
rect -3837 -381 -3747 -347
rect -3679 -381 -3589 -347
rect -3521 -381 -3431 -347
rect -3363 -381 -3273 -347
rect -3205 -381 -3115 -347
rect -3047 -381 -2957 -347
rect -2889 -381 -2799 -347
rect -2731 -381 -2641 -347
rect -2573 -381 -2483 -347
rect -2415 -381 -2325 -347
rect -2257 -381 -2167 -347
rect -2099 -381 -2009 -347
rect -1941 -381 -1851 -347
rect -1783 -381 -1693 -347
rect -1625 -381 -1535 -347
rect -1467 -381 -1377 -347
rect -1309 -381 -1219 -347
rect -1151 -381 -1061 -347
rect -993 -381 -903 -347
rect -835 -381 -745 -347
rect -677 -381 -587 -347
rect -519 -381 -429 -347
rect -361 -381 -271 -347
rect -203 -381 -113 -347
rect -45 -381 45 -347
rect 113 -381 203 -347
rect 271 -381 361 -347
rect 429 -381 519 -347
rect 587 -381 677 -347
rect 745 -381 835 -347
rect 903 -381 993 -347
rect 1061 -381 1151 -347
rect 1219 -381 1309 -347
rect 1377 -381 1467 -347
rect 1535 -381 1625 -347
rect 1693 -381 1783 -347
rect 1851 -381 1941 -347
rect 2009 -381 2099 -347
rect 2167 -381 2257 -347
rect 2325 -381 2415 -347
rect 2483 -381 2573 -347
rect 2641 -381 2731 -347
rect 2799 -381 2889 -347
rect 2957 -381 3047 -347
rect 3115 -381 3205 -347
rect 3273 -381 3363 -347
rect 3431 -381 3521 -347
rect 3589 -381 3679 -347
rect 3747 -381 3837 -347
rect 3905 -381 3995 -347
rect 4063 -381 4153 -347
rect 4221 -381 4311 -347
rect 4379 -381 4469 -347
rect 4537 -381 4627 -347
rect 4695 -381 4785 -347
rect 4853 -381 4943 -347
rect 5011 -381 5101 -347
rect 5169 -381 5259 -347
rect 5327 -381 5417 -347
rect 5485 -381 5575 -347
rect 5643 -381 5733 -347
rect 5801 -381 5891 -347
rect 5959 -381 6049 -347
rect 6117 -381 6207 -347
rect 6275 -381 6291 -347
rect -6471 -485 -6437 -423
rect 6437 -485 6471 -423
rect 6375 -519 6471 -485
<< viali >>
rect -6471 485 -6375 519
rect -6375 485 6375 519
rect -6275 347 -6207 381
rect -6117 347 -6049 381
rect -5959 347 -5891 381
rect -5801 347 -5733 381
rect -5643 347 -5575 381
rect -5485 347 -5417 381
rect -5327 347 -5259 381
rect -5169 347 -5101 381
rect -5011 347 -4943 381
rect -4853 347 -4785 381
rect -4695 347 -4627 381
rect -4537 347 -4469 381
rect -4379 347 -4311 381
rect -4221 347 -4153 381
rect -4063 347 -3995 381
rect -3905 347 -3837 381
rect -3747 347 -3679 381
rect -3589 347 -3521 381
rect -3431 347 -3363 381
rect -3273 347 -3205 381
rect -3115 347 -3047 381
rect -2957 347 -2889 381
rect -2799 347 -2731 381
rect -2641 347 -2573 381
rect -2483 347 -2415 381
rect -2325 347 -2257 381
rect -2167 347 -2099 381
rect -2009 347 -1941 381
rect -1851 347 -1783 381
rect -1693 347 -1625 381
rect -1535 347 -1467 381
rect -1377 347 -1309 381
rect -1219 347 -1151 381
rect -1061 347 -993 381
rect -903 347 -835 381
rect -745 347 -677 381
rect -587 347 -519 381
rect -429 347 -361 381
rect -271 347 -203 381
rect -113 347 -45 381
rect 45 347 113 381
rect 203 347 271 381
rect 361 347 429 381
rect 519 347 587 381
rect 677 347 745 381
rect 835 347 903 381
rect 993 347 1061 381
rect 1151 347 1219 381
rect 1309 347 1377 381
rect 1467 347 1535 381
rect 1625 347 1693 381
rect 1783 347 1851 381
rect 1941 347 2009 381
rect 2099 347 2167 381
rect 2257 347 2325 381
rect 2415 347 2483 381
rect 2573 347 2641 381
rect 2731 347 2799 381
rect 2889 347 2957 381
rect 3047 347 3115 381
rect 3205 347 3273 381
rect 3363 347 3431 381
rect 3521 347 3589 381
rect 3679 347 3747 381
rect 3837 347 3905 381
rect 3995 347 4063 381
rect 4153 347 4221 381
rect 4311 347 4379 381
rect 4469 347 4537 381
rect 4627 347 4695 381
rect 4785 347 4853 381
rect 4943 347 5011 381
rect 5101 347 5169 381
rect 5259 347 5327 381
rect 5417 347 5485 381
rect 5575 347 5643 381
rect 5733 347 5801 381
rect 5891 347 5959 381
rect 6049 347 6117 381
rect 6207 347 6275 381
rect -6337 -288 -6303 288
rect -6179 -288 -6145 288
rect -6021 -288 -5987 288
rect -5863 -288 -5829 288
rect -5705 -288 -5671 288
rect -5547 -288 -5513 288
rect -5389 -288 -5355 288
rect -5231 -288 -5197 288
rect -5073 -288 -5039 288
rect -4915 -288 -4881 288
rect -4757 -288 -4723 288
rect -4599 -288 -4565 288
rect -4441 -288 -4407 288
rect -4283 -288 -4249 288
rect -4125 -288 -4091 288
rect -3967 -288 -3933 288
rect -3809 -288 -3775 288
rect -3651 -288 -3617 288
rect -3493 -288 -3459 288
rect -3335 -288 -3301 288
rect -3177 -288 -3143 288
rect -3019 -288 -2985 288
rect -2861 -288 -2827 288
rect -2703 -288 -2669 288
rect -2545 -288 -2511 288
rect -2387 -288 -2353 288
rect -2229 -288 -2195 288
rect -2071 -288 -2037 288
rect -1913 -288 -1879 288
rect -1755 -288 -1721 288
rect -1597 -288 -1563 288
rect -1439 -288 -1405 288
rect -1281 -288 -1247 288
rect -1123 -288 -1089 288
rect -965 -288 -931 288
rect -807 -288 -773 288
rect -649 -288 -615 288
rect -491 -288 -457 288
rect -333 -288 -299 288
rect -175 -288 -141 288
rect -17 -288 17 288
rect 141 -288 175 288
rect 299 -288 333 288
rect 457 -288 491 288
rect 615 -288 649 288
rect 773 -288 807 288
rect 931 -288 965 288
rect 1089 -288 1123 288
rect 1247 -288 1281 288
rect 1405 -288 1439 288
rect 1563 -288 1597 288
rect 1721 -288 1755 288
rect 1879 -288 1913 288
rect 2037 -288 2071 288
rect 2195 -288 2229 288
rect 2353 -288 2387 288
rect 2511 -288 2545 288
rect 2669 -288 2703 288
rect 2827 -288 2861 288
rect 2985 -288 3019 288
rect 3143 -288 3177 288
rect 3301 -288 3335 288
rect 3459 -288 3493 288
rect 3617 -288 3651 288
rect 3775 -288 3809 288
rect 3933 -288 3967 288
rect 4091 -288 4125 288
rect 4249 -288 4283 288
rect 4407 -288 4441 288
rect 4565 -288 4599 288
rect 4723 -288 4757 288
rect 4881 -288 4915 288
rect 5039 -288 5073 288
rect 5197 -288 5231 288
rect 5355 -288 5389 288
rect 5513 -288 5547 288
rect 5671 -288 5705 288
rect 5829 -288 5863 288
rect 5987 -288 6021 288
rect 6145 -288 6179 288
rect 6303 -288 6337 288
rect -6275 -381 -6207 -347
rect -6117 -381 -6049 -347
rect -5959 -381 -5891 -347
rect -5801 -381 -5733 -347
rect -5643 -381 -5575 -347
rect -5485 -381 -5417 -347
rect -5327 -381 -5259 -347
rect -5169 -381 -5101 -347
rect -5011 -381 -4943 -347
rect -4853 -381 -4785 -347
rect -4695 -381 -4627 -347
rect -4537 -381 -4469 -347
rect -4379 -381 -4311 -347
rect -4221 -381 -4153 -347
rect -4063 -381 -3995 -347
rect -3905 -381 -3837 -347
rect -3747 -381 -3679 -347
rect -3589 -381 -3521 -347
rect -3431 -381 -3363 -347
rect -3273 -381 -3205 -347
rect -3115 -381 -3047 -347
rect -2957 -381 -2889 -347
rect -2799 -381 -2731 -347
rect -2641 -381 -2573 -347
rect -2483 -381 -2415 -347
rect -2325 -381 -2257 -347
rect -2167 -381 -2099 -347
rect -2009 -381 -1941 -347
rect -1851 -381 -1783 -347
rect -1693 -381 -1625 -347
rect -1535 -381 -1467 -347
rect -1377 -381 -1309 -347
rect -1219 -381 -1151 -347
rect -1061 -381 -993 -347
rect -903 -381 -835 -347
rect -745 -381 -677 -347
rect -587 -381 -519 -347
rect -429 -381 -361 -347
rect -271 -381 -203 -347
rect -113 -381 -45 -347
rect 45 -381 113 -347
rect 203 -381 271 -347
rect 361 -381 429 -347
rect 519 -381 587 -347
rect 677 -381 745 -347
rect 835 -381 903 -347
rect 993 -381 1061 -347
rect 1151 -381 1219 -347
rect 1309 -381 1377 -347
rect 1467 -381 1535 -347
rect 1625 -381 1693 -347
rect 1783 -381 1851 -347
rect 1941 -381 2009 -347
rect 2099 -381 2167 -347
rect 2257 -381 2325 -347
rect 2415 -381 2483 -347
rect 2573 -381 2641 -347
rect 2731 -381 2799 -347
rect 2889 -381 2957 -347
rect 3047 -381 3115 -347
rect 3205 -381 3273 -347
rect 3363 -381 3431 -347
rect 3521 -381 3589 -347
rect 3679 -381 3747 -347
rect 3837 -381 3905 -347
rect 3995 -381 4063 -347
rect 4153 -381 4221 -347
rect 4311 -381 4379 -347
rect 4469 -381 4537 -347
rect 4627 -381 4695 -347
rect 4785 -381 4853 -347
rect 4943 -381 5011 -347
rect 5101 -381 5169 -347
rect 5259 -381 5327 -347
rect 5417 -381 5485 -347
rect 5575 -381 5643 -347
rect 5733 -381 5801 -347
rect 5891 -381 5959 -347
rect 6049 -381 6117 -347
rect 6207 -381 6275 -347
rect 6437 -423 6471 423
rect -6471 -519 -6375 -485
rect -6375 -519 6375 -485
<< metal1 >>
rect -6483 519 6477 525
rect -6483 485 -6471 519
rect 6375 485 6477 519
rect -6483 479 6477 485
rect 6431 423 6477 479
rect -6483 381 6287 387
rect -6483 347 -6275 381
rect -6207 347 -6117 381
rect -6049 347 -5959 381
rect -5891 347 -5801 381
rect -5733 347 -5643 381
rect -5575 347 -5485 381
rect -5417 347 -5327 381
rect -5259 347 -5169 381
rect -5101 347 -5011 381
rect -4943 347 -4853 381
rect -4785 347 -4695 381
rect -4627 347 -4537 381
rect -4469 347 -4379 381
rect -4311 347 -4221 381
rect -4153 347 -4063 381
rect -3995 347 -3905 381
rect -3837 347 -3747 381
rect -3679 347 -3589 381
rect -3521 347 -3431 381
rect -3363 347 -3273 381
rect -3205 347 -3115 381
rect -3047 347 -2957 381
rect -2889 347 -2799 381
rect -2731 347 -2641 381
rect -2573 347 -2483 381
rect -2415 347 -2325 381
rect -2257 347 -2167 381
rect -2099 347 -2009 381
rect -1941 347 -1851 381
rect -1783 347 -1693 381
rect -1625 347 -1535 381
rect -1467 347 -1377 381
rect -1309 347 -1219 381
rect -1151 347 -1061 381
rect -993 347 -903 381
rect -835 347 -745 381
rect -677 347 -587 381
rect -519 347 -429 381
rect -361 347 -271 381
rect -203 347 -113 381
rect -45 347 45 381
rect 113 347 203 381
rect 271 347 361 381
rect 429 347 519 381
rect 587 347 677 381
rect 745 347 835 381
rect 903 347 993 381
rect 1061 347 1151 381
rect 1219 347 1309 381
rect 1377 347 1467 381
rect 1535 347 1625 381
rect 1693 347 1783 381
rect 1851 347 1941 381
rect 2009 347 2099 381
rect 2167 347 2257 381
rect 2325 347 2415 381
rect 2483 347 2573 381
rect 2641 347 2731 381
rect 2799 347 2889 381
rect 2957 347 3047 381
rect 3115 347 3205 381
rect 3273 347 3363 381
rect 3431 347 3521 381
rect 3589 347 3679 381
rect 3747 347 3837 381
rect 3905 347 3995 381
rect 4063 347 4153 381
rect 4221 347 4311 381
rect 4379 347 4469 381
rect 4537 347 4627 381
rect 4695 347 4785 381
rect 4853 347 4943 381
rect 5011 347 5101 381
rect 5169 347 5259 381
rect 5327 347 5417 381
rect 5485 347 5575 381
rect 5643 347 5733 381
rect 5801 347 5891 381
rect 5959 347 6049 381
rect 6117 347 6207 381
rect 6275 347 6287 381
rect -6483 341 6287 347
rect -6483 -341 -6437 341
rect -6346 288 -6294 300
rect -6346 -26 -6337 288
rect -6303 -26 -6294 288
rect -6346 -300 -6294 -294
rect -6188 294 -6136 300
rect -6188 -288 -6179 26
rect -6145 -288 -6136 26
rect -6188 -300 -6136 -288
rect -6030 288 -5978 300
rect -6030 -26 -6021 288
rect -5987 -26 -5978 288
rect -6030 -300 -5978 -294
rect -5872 294 -5820 300
rect -5872 -288 -5863 26
rect -5829 -288 -5820 26
rect -5872 -300 -5820 -288
rect -5714 288 -5662 300
rect -5714 -26 -5705 288
rect -5671 -26 -5662 288
rect -5714 -300 -5662 -294
rect -5556 294 -5504 300
rect -5556 -288 -5547 26
rect -5513 -288 -5504 26
rect -5556 -300 -5504 -288
rect -5398 288 -5346 300
rect -5398 -26 -5389 288
rect -5355 -26 -5346 288
rect -5398 -300 -5346 -294
rect -5240 294 -5188 300
rect -5240 -288 -5231 26
rect -5197 -288 -5188 26
rect -5240 -300 -5188 -288
rect -5082 288 -5030 300
rect -5082 -26 -5073 288
rect -5039 -26 -5030 288
rect -5082 -300 -5030 -294
rect -4924 294 -4872 300
rect -4924 -288 -4915 26
rect -4881 -288 -4872 26
rect -4924 -300 -4872 -288
rect -4766 288 -4714 300
rect -4766 -26 -4757 288
rect -4723 -26 -4714 288
rect -4766 -300 -4714 -294
rect -4608 294 -4556 300
rect -4608 -288 -4599 26
rect -4565 -288 -4556 26
rect -4608 -300 -4556 -288
rect -4450 288 -4398 300
rect -4450 -26 -4441 288
rect -4407 -26 -4398 288
rect -4450 -300 -4398 -294
rect -4292 294 -4240 300
rect -4292 -288 -4283 26
rect -4249 -288 -4240 26
rect -4292 -300 -4240 -288
rect -4134 288 -4082 300
rect -4134 -26 -4125 288
rect -4091 -26 -4082 288
rect -4134 -300 -4082 -294
rect -3976 294 -3924 300
rect -3976 -288 -3967 26
rect -3933 -288 -3924 26
rect -3976 -300 -3924 -288
rect -3818 288 -3766 300
rect -3818 -26 -3809 288
rect -3775 -26 -3766 288
rect -3818 -300 -3766 -294
rect -3660 294 -3608 300
rect -3660 -288 -3651 26
rect -3617 -288 -3608 26
rect -3660 -300 -3608 -288
rect -3502 288 -3450 300
rect -3502 -26 -3493 288
rect -3459 -26 -3450 288
rect -3502 -300 -3450 -294
rect -3344 294 -3292 300
rect -3344 -288 -3335 26
rect -3301 -288 -3292 26
rect -3344 -300 -3292 -288
rect -3186 288 -3134 300
rect -3186 -26 -3177 288
rect -3143 -26 -3134 288
rect -3186 -300 -3134 -294
rect -3028 294 -2976 300
rect -3028 -288 -3019 26
rect -2985 -288 -2976 26
rect -3028 -300 -2976 -288
rect -2870 288 -2818 300
rect -2870 -26 -2861 288
rect -2827 -26 -2818 288
rect -2870 -300 -2818 -294
rect -2712 294 -2660 300
rect -2712 -288 -2703 26
rect -2669 -288 -2660 26
rect -2712 -300 -2660 -288
rect -2554 288 -2502 300
rect -2554 -26 -2545 288
rect -2511 -26 -2502 288
rect -2554 -300 -2502 -294
rect -2396 294 -2344 300
rect -2396 -288 -2387 26
rect -2353 -288 -2344 26
rect -2396 -300 -2344 -288
rect -2238 288 -2186 300
rect -2238 -26 -2229 288
rect -2195 -26 -2186 288
rect -2238 -300 -2186 -294
rect -2080 294 -2028 300
rect -2080 -288 -2071 26
rect -2037 -288 -2028 26
rect -2080 -300 -2028 -288
rect -1922 288 -1870 300
rect -1922 -26 -1913 288
rect -1879 -26 -1870 288
rect -1922 -300 -1870 -294
rect -1764 294 -1712 300
rect -1764 -288 -1755 26
rect -1721 -288 -1712 26
rect -1764 -300 -1712 -288
rect -1606 288 -1554 300
rect -1606 -26 -1597 288
rect -1563 -26 -1554 288
rect -1606 -300 -1554 -294
rect -1448 294 -1396 300
rect -1448 -288 -1439 26
rect -1405 -288 -1396 26
rect -1448 -300 -1396 -288
rect -1290 288 -1238 300
rect -1290 -26 -1281 288
rect -1247 -26 -1238 288
rect -1290 -300 -1238 -294
rect -1132 294 -1080 300
rect -1132 -288 -1123 26
rect -1089 -288 -1080 26
rect -1132 -300 -1080 -288
rect -974 288 -922 300
rect -974 -26 -965 288
rect -931 -26 -922 288
rect -974 -300 -922 -294
rect -816 294 -764 300
rect -816 -288 -807 26
rect -773 -288 -764 26
rect -816 -300 -764 -288
rect -658 288 -606 300
rect -658 -26 -649 288
rect -615 -26 -606 288
rect -658 -300 -606 -294
rect -500 294 -448 300
rect -500 -288 -491 26
rect -457 -288 -448 26
rect -500 -300 -448 -288
rect -342 288 -290 300
rect -342 -26 -333 288
rect -299 -26 -290 288
rect -342 -300 -290 -294
rect -184 294 -132 300
rect -184 -288 -175 26
rect -141 -288 -132 26
rect -184 -300 -132 -288
rect -26 288 26 300
rect -26 -26 -17 288
rect 17 -26 26 288
rect -26 -300 26 -294
rect 132 294 184 300
rect 132 -288 141 26
rect 175 -288 184 26
rect 132 -300 184 -288
rect 290 288 342 300
rect 290 -26 299 288
rect 333 -26 342 288
rect 290 -300 342 -294
rect 448 294 500 300
rect 448 -288 457 26
rect 491 -288 500 26
rect 448 -300 500 -288
rect 606 288 658 300
rect 606 -26 615 288
rect 649 -26 658 288
rect 606 -300 658 -294
rect 764 294 816 300
rect 764 -288 773 26
rect 807 -288 816 26
rect 764 -300 816 -288
rect 922 288 974 300
rect 922 -26 931 288
rect 965 -26 974 288
rect 922 -300 974 -294
rect 1080 294 1132 300
rect 1080 -288 1089 26
rect 1123 -288 1132 26
rect 1080 -300 1132 -288
rect 1238 288 1290 300
rect 1238 -26 1247 288
rect 1281 -26 1290 288
rect 1238 -300 1290 -294
rect 1396 294 1448 300
rect 1396 -288 1405 26
rect 1439 -288 1448 26
rect 1396 -300 1448 -288
rect 1554 288 1606 300
rect 1554 -26 1563 288
rect 1597 -26 1606 288
rect 1554 -300 1606 -294
rect 1712 294 1764 300
rect 1712 -288 1721 26
rect 1755 -288 1764 26
rect 1712 -300 1764 -288
rect 1870 288 1922 300
rect 1870 -26 1879 288
rect 1913 -26 1922 288
rect 1870 -300 1922 -294
rect 2028 294 2080 300
rect 2028 -288 2037 26
rect 2071 -288 2080 26
rect 2028 -300 2080 -288
rect 2186 288 2238 300
rect 2186 -26 2195 288
rect 2229 -26 2238 288
rect 2186 -300 2238 -294
rect 2344 294 2396 300
rect 2344 -288 2353 26
rect 2387 -288 2396 26
rect 2344 -300 2396 -288
rect 2502 288 2554 300
rect 2502 -26 2511 288
rect 2545 -26 2554 288
rect 2502 -300 2554 -294
rect 2660 294 2712 300
rect 2660 -288 2669 26
rect 2703 -288 2712 26
rect 2660 -300 2712 -288
rect 2818 288 2870 300
rect 2818 -26 2827 288
rect 2861 -26 2870 288
rect 2818 -300 2870 -294
rect 2976 294 3028 300
rect 2976 -288 2985 26
rect 3019 -288 3028 26
rect 2976 -300 3028 -288
rect 3134 288 3186 300
rect 3134 -26 3143 288
rect 3177 -26 3186 288
rect 3134 -300 3186 -294
rect 3292 294 3344 300
rect 3292 -288 3301 26
rect 3335 -288 3344 26
rect 3292 -300 3344 -288
rect 3450 288 3502 300
rect 3450 -26 3459 288
rect 3493 -26 3502 288
rect 3450 -300 3502 -294
rect 3608 294 3660 300
rect 3608 -288 3617 26
rect 3651 -288 3660 26
rect 3608 -300 3660 -288
rect 3766 288 3818 300
rect 3766 -26 3775 288
rect 3809 -26 3818 288
rect 3766 -300 3818 -294
rect 3924 294 3976 300
rect 3924 -288 3933 26
rect 3967 -288 3976 26
rect 3924 -300 3976 -288
rect 4082 288 4134 300
rect 4082 -26 4091 288
rect 4125 -26 4134 288
rect 4082 -300 4134 -294
rect 4240 294 4292 300
rect 4240 -288 4249 26
rect 4283 -288 4292 26
rect 4240 -300 4292 -288
rect 4398 288 4450 300
rect 4398 -26 4407 288
rect 4441 -26 4450 288
rect 4398 -300 4450 -294
rect 4556 294 4608 300
rect 4556 -288 4565 26
rect 4599 -288 4608 26
rect 4556 -300 4608 -288
rect 4714 288 4766 300
rect 4714 -26 4723 288
rect 4757 -26 4766 288
rect 4714 -300 4766 -294
rect 4872 294 4924 300
rect 4872 -288 4881 26
rect 4915 -288 4924 26
rect 4872 -300 4924 -288
rect 5030 288 5082 300
rect 5030 -26 5039 288
rect 5073 -26 5082 288
rect 5030 -300 5082 -294
rect 5188 294 5240 300
rect 5188 -288 5197 26
rect 5231 -288 5240 26
rect 5188 -300 5240 -288
rect 5346 288 5398 300
rect 5346 -26 5355 288
rect 5389 -26 5398 288
rect 5346 -300 5398 -294
rect 5504 294 5556 300
rect 5504 -288 5513 26
rect 5547 -288 5556 26
rect 5504 -300 5556 -288
rect 5662 288 5714 300
rect 5662 -26 5671 288
rect 5705 -26 5714 288
rect 5662 -300 5714 -294
rect 5820 294 5872 300
rect 5820 -288 5829 26
rect 5863 -288 5872 26
rect 5820 -300 5872 -288
rect 5978 288 6030 300
rect 5978 -26 5987 288
rect 6021 -26 6030 288
rect 5978 -300 6030 -294
rect 6136 294 6188 300
rect 6136 -288 6145 26
rect 6179 -288 6188 26
rect 6136 -300 6188 -288
rect 6294 288 6346 300
rect 6294 -26 6303 288
rect 6337 -26 6346 288
rect 6294 -300 6346 -294
rect -6483 -347 6287 -341
rect -6483 -381 -6275 -347
rect -6207 -381 -6117 -347
rect -6049 -381 -5959 -347
rect -5891 -381 -5801 -347
rect -5733 -381 -5643 -347
rect -5575 -381 -5485 -347
rect -5417 -381 -5327 -347
rect -5259 -381 -5169 -347
rect -5101 -381 -5011 -347
rect -4943 -381 -4853 -347
rect -4785 -381 -4695 -347
rect -4627 -381 -4537 -347
rect -4469 -381 -4379 -347
rect -4311 -381 -4221 -347
rect -4153 -381 -4063 -347
rect -3995 -381 -3905 -347
rect -3837 -381 -3747 -347
rect -3679 -381 -3589 -347
rect -3521 -381 -3431 -347
rect -3363 -381 -3273 -347
rect -3205 -381 -3115 -347
rect -3047 -381 -2957 -347
rect -2889 -381 -2799 -347
rect -2731 -381 -2641 -347
rect -2573 -381 -2483 -347
rect -2415 -381 -2325 -347
rect -2257 -381 -2167 -347
rect -2099 -381 -2009 -347
rect -1941 -381 -1851 -347
rect -1783 -381 -1693 -347
rect -1625 -381 -1535 -347
rect -1467 -381 -1377 -347
rect -1309 -381 -1219 -347
rect -1151 -381 -1061 -347
rect -993 -381 -903 -347
rect -835 -381 -745 -347
rect -677 -381 -587 -347
rect -519 -381 -429 -347
rect -361 -381 -271 -347
rect -203 -381 -113 -347
rect -45 -381 45 -347
rect 113 -381 203 -347
rect 271 -381 361 -347
rect 429 -381 519 -347
rect 587 -381 677 -347
rect 745 -381 835 -347
rect 903 -381 993 -347
rect 1061 -381 1151 -347
rect 1219 -381 1309 -347
rect 1377 -381 1467 -347
rect 1535 -381 1625 -347
rect 1693 -381 1783 -347
rect 1851 -381 1941 -347
rect 2009 -381 2099 -347
rect 2167 -381 2257 -347
rect 2325 -381 2415 -347
rect 2483 -381 2573 -347
rect 2641 -381 2731 -347
rect 2799 -381 2889 -347
rect 2957 -381 3047 -347
rect 3115 -381 3205 -347
rect 3273 -381 3363 -347
rect 3431 -381 3521 -347
rect 3589 -381 3679 -347
rect 3747 -381 3837 -347
rect 3905 -381 3995 -347
rect 4063 -381 4153 -347
rect 4221 -381 4311 -347
rect 4379 -381 4469 -347
rect 4537 -381 4627 -347
rect 4695 -381 4785 -347
rect 4853 -381 4943 -347
rect 5011 -381 5101 -347
rect 5169 -381 5259 -347
rect 5327 -381 5417 -347
rect 5485 -381 5575 -347
rect 5643 -381 5733 -347
rect 5801 -381 5891 -347
rect 5959 -381 6049 -347
rect 6117 -381 6207 -347
rect 6275 -381 6287 -347
rect -6483 -387 6287 -381
rect 6431 -423 6437 423
rect 6471 -423 6477 423
rect 6431 -479 6477 -423
rect -6483 -485 6477 -479
rect -6483 -519 -6471 -485
rect 6375 -519 6477 -485
rect -6483 -525 6477 -519
<< via1 >>
rect -6346 -288 -6337 -26
rect -6337 -288 -6303 -26
rect -6303 -288 -6294 -26
rect -6346 -294 -6294 -288
rect -6188 288 -6136 294
rect -6188 26 -6179 288
rect -6179 26 -6145 288
rect -6145 26 -6136 288
rect -6030 -288 -6021 -26
rect -6021 -288 -5987 -26
rect -5987 -288 -5978 -26
rect -6030 -294 -5978 -288
rect -5872 288 -5820 294
rect -5872 26 -5863 288
rect -5863 26 -5829 288
rect -5829 26 -5820 288
rect -5714 -288 -5705 -26
rect -5705 -288 -5671 -26
rect -5671 -288 -5662 -26
rect -5714 -294 -5662 -288
rect -5556 288 -5504 294
rect -5556 26 -5547 288
rect -5547 26 -5513 288
rect -5513 26 -5504 288
rect -5398 -288 -5389 -26
rect -5389 -288 -5355 -26
rect -5355 -288 -5346 -26
rect -5398 -294 -5346 -288
rect -5240 288 -5188 294
rect -5240 26 -5231 288
rect -5231 26 -5197 288
rect -5197 26 -5188 288
rect -5082 -288 -5073 -26
rect -5073 -288 -5039 -26
rect -5039 -288 -5030 -26
rect -5082 -294 -5030 -288
rect -4924 288 -4872 294
rect -4924 26 -4915 288
rect -4915 26 -4881 288
rect -4881 26 -4872 288
rect -4766 -288 -4757 -26
rect -4757 -288 -4723 -26
rect -4723 -288 -4714 -26
rect -4766 -294 -4714 -288
rect -4608 288 -4556 294
rect -4608 26 -4599 288
rect -4599 26 -4565 288
rect -4565 26 -4556 288
rect -4450 -288 -4441 -26
rect -4441 -288 -4407 -26
rect -4407 -288 -4398 -26
rect -4450 -294 -4398 -288
rect -4292 288 -4240 294
rect -4292 26 -4283 288
rect -4283 26 -4249 288
rect -4249 26 -4240 288
rect -4134 -288 -4125 -26
rect -4125 -288 -4091 -26
rect -4091 -288 -4082 -26
rect -4134 -294 -4082 -288
rect -3976 288 -3924 294
rect -3976 26 -3967 288
rect -3967 26 -3933 288
rect -3933 26 -3924 288
rect -3818 -288 -3809 -26
rect -3809 -288 -3775 -26
rect -3775 -288 -3766 -26
rect -3818 -294 -3766 -288
rect -3660 288 -3608 294
rect -3660 26 -3651 288
rect -3651 26 -3617 288
rect -3617 26 -3608 288
rect -3502 -288 -3493 -26
rect -3493 -288 -3459 -26
rect -3459 -288 -3450 -26
rect -3502 -294 -3450 -288
rect -3344 288 -3292 294
rect -3344 26 -3335 288
rect -3335 26 -3301 288
rect -3301 26 -3292 288
rect -3186 -288 -3177 -26
rect -3177 -288 -3143 -26
rect -3143 -288 -3134 -26
rect -3186 -294 -3134 -288
rect -3028 288 -2976 294
rect -3028 26 -3019 288
rect -3019 26 -2985 288
rect -2985 26 -2976 288
rect -2870 -288 -2861 -26
rect -2861 -288 -2827 -26
rect -2827 -288 -2818 -26
rect -2870 -294 -2818 -288
rect -2712 288 -2660 294
rect -2712 26 -2703 288
rect -2703 26 -2669 288
rect -2669 26 -2660 288
rect -2554 -288 -2545 -26
rect -2545 -288 -2511 -26
rect -2511 -288 -2502 -26
rect -2554 -294 -2502 -288
rect -2396 288 -2344 294
rect -2396 26 -2387 288
rect -2387 26 -2353 288
rect -2353 26 -2344 288
rect -2238 -288 -2229 -26
rect -2229 -288 -2195 -26
rect -2195 -288 -2186 -26
rect -2238 -294 -2186 -288
rect -2080 288 -2028 294
rect -2080 26 -2071 288
rect -2071 26 -2037 288
rect -2037 26 -2028 288
rect -1922 -288 -1913 -26
rect -1913 -288 -1879 -26
rect -1879 -288 -1870 -26
rect -1922 -294 -1870 -288
rect -1764 288 -1712 294
rect -1764 26 -1755 288
rect -1755 26 -1721 288
rect -1721 26 -1712 288
rect -1606 -288 -1597 -26
rect -1597 -288 -1563 -26
rect -1563 -288 -1554 -26
rect -1606 -294 -1554 -288
rect -1448 288 -1396 294
rect -1448 26 -1439 288
rect -1439 26 -1405 288
rect -1405 26 -1396 288
rect -1290 -288 -1281 -26
rect -1281 -288 -1247 -26
rect -1247 -288 -1238 -26
rect -1290 -294 -1238 -288
rect -1132 288 -1080 294
rect -1132 26 -1123 288
rect -1123 26 -1089 288
rect -1089 26 -1080 288
rect -974 -288 -965 -26
rect -965 -288 -931 -26
rect -931 -288 -922 -26
rect -974 -294 -922 -288
rect -816 288 -764 294
rect -816 26 -807 288
rect -807 26 -773 288
rect -773 26 -764 288
rect -658 -288 -649 -26
rect -649 -288 -615 -26
rect -615 -288 -606 -26
rect -658 -294 -606 -288
rect -500 288 -448 294
rect -500 26 -491 288
rect -491 26 -457 288
rect -457 26 -448 288
rect -342 -288 -333 -26
rect -333 -288 -299 -26
rect -299 -288 -290 -26
rect -342 -294 -290 -288
rect -184 288 -132 294
rect -184 26 -175 288
rect -175 26 -141 288
rect -141 26 -132 288
rect -26 -288 -17 -26
rect -17 -288 17 -26
rect 17 -288 26 -26
rect -26 -294 26 -288
rect 132 288 184 294
rect 132 26 141 288
rect 141 26 175 288
rect 175 26 184 288
rect 290 -288 299 -26
rect 299 -288 333 -26
rect 333 -288 342 -26
rect 290 -294 342 -288
rect 448 288 500 294
rect 448 26 457 288
rect 457 26 491 288
rect 491 26 500 288
rect 606 -288 615 -26
rect 615 -288 649 -26
rect 649 -288 658 -26
rect 606 -294 658 -288
rect 764 288 816 294
rect 764 26 773 288
rect 773 26 807 288
rect 807 26 816 288
rect 922 -288 931 -26
rect 931 -288 965 -26
rect 965 -288 974 -26
rect 922 -294 974 -288
rect 1080 288 1132 294
rect 1080 26 1089 288
rect 1089 26 1123 288
rect 1123 26 1132 288
rect 1238 -288 1247 -26
rect 1247 -288 1281 -26
rect 1281 -288 1290 -26
rect 1238 -294 1290 -288
rect 1396 288 1448 294
rect 1396 26 1405 288
rect 1405 26 1439 288
rect 1439 26 1448 288
rect 1554 -288 1563 -26
rect 1563 -288 1597 -26
rect 1597 -288 1606 -26
rect 1554 -294 1606 -288
rect 1712 288 1764 294
rect 1712 26 1721 288
rect 1721 26 1755 288
rect 1755 26 1764 288
rect 1870 -288 1879 -26
rect 1879 -288 1913 -26
rect 1913 -288 1922 -26
rect 1870 -294 1922 -288
rect 2028 288 2080 294
rect 2028 26 2037 288
rect 2037 26 2071 288
rect 2071 26 2080 288
rect 2186 -288 2195 -26
rect 2195 -288 2229 -26
rect 2229 -288 2238 -26
rect 2186 -294 2238 -288
rect 2344 288 2396 294
rect 2344 26 2353 288
rect 2353 26 2387 288
rect 2387 26 2396 288
rect 2502 -288 2511 -26
rect 2511 -288 2545 -26
rect 2545 -288 2554 -26
rect 2502 -294 2554 -288
rect 2660 288 2712 294
rect 2660 26 2669 288
rect 2669 26 2703 288
rect 2703 26 2712 288
rect 2818 -288 2827 -26
rect 2827 -288 2861 -26
rect 2861 -288 2870 -26
rect 2818 -294 2870 -288
rect 2976 288 3028 294
rect 2976 26 2985 288
rect 2985 26 3019 288
rect 3019 26 3028 288
rect 3134 -288 3143 -26
rect 3143 -288 3177 -26
rect 3177 -288 3186 -26
rect 3134 -294 3186 -288
rect 3292 288 3344 294
rect 3292 26 3301 288
rect 3301 26 3335 288
rect 3335 26 3344 288
rect 3450 -288 3459 -26
rect 3459 -288 3493 -26
rect 3493 -288 3502 -26
rect 3450 -294 3502 -288
rect 3608 288 3660 294
rect 3608 26 3617 288
rect 3617 26 3651 288
rect 3651 26 3660 288
rect 3766 -288 3775 -26
rect 3775 -288 3809 -26
rect 3809 -288 3818 -26
rect 3766 -294 3818 -288
rect 3924 288 3976 294
rect 3924 26 3933 288
rect 3933 26 3967 288
rect 3967 26 3976 288
rect 4082 -288 4091 -26
rect 4091 -288 4125 -26
rect 4125 -288 4134 -26
rect 4082 -294 4134 -288
rect 4240 288 4292 294
rect 4240 26 4249 288
rect 4249 26 4283 288
rect 4283 26 4292 288
rect 4398 -288 4407 -26
rect 4407 -288 4441 -26
rect 4441 -288 4450 -26
rect 4398 -294 4450 -288
rect 4556 288 4608 294
rect 4556 26 4565 288
rect 4565 26 4599 288
rect 4599 26 4608 288
rect 4714 -288 4723 -26
rect 4723 -288 4757 -26
rect 4757 -288 4766 -26
rect 4714 -294 4766 -288
rect 4872 288 4924 294
rect 4872 26 4881 288
rect 4881 26 4915 288
rect 4915 26 4924 288
rect 5030 -288 5039 -26
rect 5039 -288 5073 -26
rect 5073 -288 5082 -26
rect 5030 -294 5082 -288
rect 5188 288 5240 294
rect 5188 26 5197 288
rect 5197 26 5231 288
rect 5231 26 5240 288
rect 5346 -288 5355 -26
rect 5355 -288 5389 -26
rect 5389 -288 5398 -26
rect 5346 -294 5398 -288
rect 5504 288 5556 294
rect 5504 26 5513 288
rect 5513 26 5547 288
rect 5547 26 5556 288
rect 5662 -288 5671 -26
rect 5671 -288 5705 -26
rect 5705 -288 5714 -26
rect 5662 -294 5714 -288
rect 5820 288 5872 294
rect 5820 26 5829 288
rect 5829 26 5863 288
rect 5863 26 5872 288
rect 5978 -288 5987 -26
rect 5987 -288 6021 -26
rect 6021 -288 6030 -26
rect 5978 -294 6030 -288
rect 6136 288 6188 294
rect 6136 26 6145 288
rect 6145 26 6179 288
rect 6179 26 6188 288
rect 6294 -288 6303 -26
rect 6303 -288 6337 -26
rect 6337 -288 6346 -26
rect 6294 -294 6346 -288
<< metal2 >>
rect -6188 294 6188 300
rect -6136 26 -5872 294
rect -5820 26 -5556 294
rect -5504 26 -5240 294
rect -5188 26 -4924 294
rect -4872 26 -4608 294
rect -4556 26 -4292 294
rect -4240 26 -3976 294
rect -3924 26 -3660 294
rect -3608 26 -3344 294
rect -3292 26 -3028 294
rect -2976 26 -2712 294
rect -2660 26 -2396 294
rect -2344 26 -2080 294
rect -2028 26 -1764 294
rect -1712 26 -1448 294
rect -1396 26 -1132 294
rect -1080 26 -816 294
rect -764 26 -500 294
rect -448 26 -184 294
rect -132 26 132 294
rect 184 26 448 294
rect 500 26 764 294
rect 816 26 1080 294
rect 1132 26 1396 294
rect 1448 26 1712 294
rect 1764 26 2028 294
rect 2080 26 2344 294
rect 2396 26 2660 294
rect 2712 26 2976 294
rect 3028 26 3292 294
rect 3344 26 3608 294
rect 3660 26 3924 294
rect 3976 26 4240 294
rect 4292 26 4556 294
rect 4608 26 4872 294
rect 4924 26 5188 294
rect 5240 26 5504 294
rect 5556 26 5820 294
rect 5872 26 6136 294
rect -6188 20 6188 26
rect -6346 -26 6346 -20
rect -6294 -294 -6030 -26
rect -5978 -294 -5714 -26
rect -5662 -294 -5398 -26
rect -5346 -294 -5082 -26
rect -5030 -294 -4766 -26
rect -4714 -294 -4450 -26
rect -4398 -294 -4134 -26
rect -4082 -294 -3818 -26
rect -3766 -294 -3502 -26
rect -3450 -294 -3186 -26
rect -3134 -294 -2870 -26
rect -2818 -294 -2554 -26
rect -2502 -294 -2238 -26
rect -2186 -294 -1922 -26
rect -1870 -294 -1606 -26
rect -1554 -294 -1290 -26
rect -1238 -294 -974 -26
rect -922 -294 -658 -26
rect -606 -294 -342 -26
rect -290 -294 -26 -26
rect 26 -294 290 -26
rect 342 -294 606 -26
rect 658 -294 922 -26
rect 974 -294 1238 -26
rect 1290 -294 1554 -26
rect 1606 -294 1870 -26
rect 1922 -294 2186 -26
rect 2238 -294 2502 -26
rect 2554 -294 2818 -26
rect 2870 -294 3134 -26
rect 3186 -294 3450 -26
rect 3502 -294 3766 -26
rect 3818 -294 4082 -26
rect 4134 -294 4398 -26
rect 4450 -294 4714 -26
rect 4766 -294 5030 -26
rect 5082 -294 5346 -26
rect 5398 -294 5662 -26
rect 5714 -294 5978 -26
rect 6030 -294 6294 -26
rect -6346 -300 6346 -294
<< properties >>
string FIXED_BBOX -6454 -502 6454 502
string gencell sky130_fd_pr__pfet_g5v0d10v5
string library sky130
string parameters w 3 l 0.5 m 1 nf 80 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
