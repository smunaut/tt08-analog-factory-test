magic
tech sky130A
magscale 1 2
timestamp 1725098041
<< pwell >>
rect -13155 -658 13155 658
<< mvnmos >>
rect -12927 -400 -12827 400
rect -12769 -400 -12669 400
rect -12611 -400 -12511 400
rect -12453 -400 -12353 400
rect -12295 -400 -12195 400
rect -12137 -400 -12037 400
rect -11979 -400 -11879 400
rect -11821 -400 -11721 400
rect -11663 -400 -11563 400
rect -11505 -400 -11405 400
rect -11347 -400 -11247 400
rect -11189 -400 -11089 400
rect -11031 -400 -10931 400
rect -10873 -400 -10773 400
rect -10715 -400 -10615 400
rect -10557 -400 -10457 400
rect -10399 -400 -10299 400
rect -10241 -400 -10141 400
rect -10083 -400 -9983 400
rect -9925 -400 -9825 400
rect -9767 -400 -9667 400
rect -9609 -400 -9509 400
rect -9451 -400 -9351 400
rect -9293 -400 -9193 400
rect -9135 -400 -9035 400
rect -8977 -400 -8877 400
rect -8819 -400 -8719 400
rect -8661 -400 -8561 400
rect -8503 -400 -8403 400
rect -8345 -400 -8245 400
rect -8187 -400 -8087 400
rect -8029 -400 -7929 400
rect -7871 -400 -7771 400
rect -7713 -400 -7613 400
rect -7555 -400 -7455 400
rect -7397 -400 -7297 400
rect -7239 -400 -7139 400
rect -7081 -400 -6981 400
rect -6923 -400 -6823 400
rect -6765 -400 -6665 400
rect -6607 -400 -6507 400
rect -6449 -400 -6349 400
rect -6291 -400 -6191 400
rect -6133 -400 -6033 400
rect -5975 -400 -5875 400
rect -5817 -400 -5717 400
rect -5659 -400 -5559 400
rect -5501 -400 -5401 400
rect -5343 -400 -5243 400
rect -5185 -400 -5085 400
rect -5027 -400 -4927 400
rect -4869 -400 -4769 400
rect -4711 -400 -4611 400
rect -4553 -400 -4453 400
rect -4395 -400 -4295 400
rect -4237 -400 -4137 400
rect -4079 -400 -3979 400
rect -3921 -400 -3821 400
rect -3763 -400 -3663 400
rect -3605 -400 -3505 400
rect -3447 -400 -3347 400
rect -3289 -400 -3189 400
rect -3131 -400 -3031 400
rect -2973 -400 -2873 400
rect -2815 -400 -2715 400
rect -2657 -400 -2557 400
rect -2499 -400 -2399 400
rect -2341 -400 -2241 400
rect -2183 -400 -2083 400
rect -2025 -400 -1925 400
rect -1867 -400 -1767 400
rect -1709 -400 -1609 400
rect -1551 -400 -1451 400
rect -1393 -400 -1293 400
rect -1235 -400 -1135 400
rect -1077 -400 -977 400
rect -919 -400 -819 400
rect -761 -400 -661 400
rect -603 -400 -503 400
rect -445 -400 -345 400
rect -287 -400 -187 400
rect -129 -400 -29 400
rect 29 -400 129 400
rect 187 -400 287 400
rect 345 -400 445 400
rect 503 -400 603 400
rect 661 -400 761 400
rect 819 -400 919 400
rect 977 -400 1077 400
rect 1135 -400 1235 400
rect 1293 -400 1393 400
rect 1451 -400 1551 400
rect 1609 -400 1709 400
rect 1767 -400 1867 400
rect 1925 -400 2025 400
rect 2083 -400 2183 400
rect 2241 -400 2341 400
rect 2399 -400 2499 400
rect 2557 -400 2657 400
rect 2715 -400 2815 400
rect 2873 -400 2973 400
rect 3031 -400 3131 400
rect 3189 -400 3289 400
rect 3347 -400 3447 400
rect 3505 -400 3605 400
rect 3663 -400 3763 400
rect 3821 -400 3921 400
rect 3979 -400 4079 400
rect 4137 -400 4237 400
rect 4295 -400 4395 400
rect 4453 -400 4553 400
rect 4611 -400 4711 400
rect 4769 -400 4869 400
rect 4927 -400 5027 400
rect 5085 -400 5185 400
rect 5243 -400 5343 400
rect 5401 -400 5501 400
rect 5559 -400 5659 400
rect 5717 -400 5817 400
rect 5875 -400 5975 400
rect 6033 -400 6133 400
rect 6191 -400 6291 400
rect 6349 -400 6449 400
rect 6507 -400 6607 400
rect 6665 -400 6765 400
rect 6823 -400 6923 400
rect 6981 -400 7081 400
rect 7139 -400 7239 400
rect 7297 -400 7397 400
rect 7455 -400 7555 400
rect 7613 -400 7713 400
rect 7771 -400 7871 400
rect 7929 -400 8029 400
rect 8087 -400 8187 400
rect 8245 -400 8345 400
rect 8403 -400 8503 400
rect 8561 -400 8661 400
rect 8719 -400 8819 400
rect 8877 -400 8977 400
rect 9035 -400 9135 400
rect 9193 -400 9293 400
rect 9351 -400 9451 400
rect 9509 -400 9609 400
rect 9667 -400 9767 400
rect 9825 -400 9925 400
rect 9983 -400 10083 400
rect 10141 -400 10241 400
rect 10299 -400 10399 400
rect 10457 -400 10557 400
rect 10615 -400 10715 400
rect 10773 -400 10873 400
rect 10931 -400 11031 400
rect 11089 -400 11189 400
rect 11247 -400 11347 400
rect 11405 -400 11505 400
rect 11563 -400 11663 400
rect 11721 -400 11821 400
rect 11879 -400 11979 400
rect 12037 -400 12137 400
rect 12195 -400 12295 400
rect 12353 -400 12453 400
rect 12511 -400 12611 400
rect 12669 -400 12769 400
rect 12827 -400 12927 400
<< mvndiff >>
rect -12985 388 -12927 400
rect -12985 -388 -12973 388
rect -12939 -388 -12927 388
rect -12985 -400 -12927 -388
rect -12827 388 -12769 400
rect -12827 -388 -12815 388
rect -12781 -388 -12769 388
rect -12827 -400 -12769 -388
rect -12669 388 -12611 400
rect -12669 -388 -12657 388
rect -12623 -388 -12611 388
rect -12669 -400 -12611 -388
rect -12511 388 -12453 400
rect -12511 -388 -12499 388
rect -12465 -388 -12453 388
rect -12511 -400 -12453 -388
rect -12353 388 -12295 400
rect -12353 -388 -12341 388
rect -12307 -388 -12295 388
rect -12353 -400 -12295 -388
rect -12195 388 -12137 400
rect -12195 -388 -12183 388
rect -12149 -388 -12137 388
rect -12195 -400 -12137 -388
rect -12037 388 -11979 400
rect -12037 -388 -12025 388
rect -11991 -388 -11979 388
rect -12037 -400 -11979 -388
rect -11879 388 -11821 400
rect -11879 -388 -11867 388
rect -11833 -388 -11821 388
rect -11879 -400 -11821 -388
rect -11721 388 -11663 400
rect -11721 -388 -11709 388
rect -11675 -388 -11663 388
rect -11721 -400 -11663 -388
rect -11563 388 -11505 400
rect -11563 -388 -11551 388
rect -11517 -388 -11505 388
rect -11563 -400 -11505 -388
rect -11405 388 -11347 400
rect -11405 -388 -11393 388
rect -11359 -388 -11347 388
rect -11405 -400 -11347 -388
rect -11247 388 -11189 400
rect -11247 -388 -11235 388
rect -11201 -388 -11189 388
rect -11247 -400 -11189 -388
rect -11089 388 -11031 400
rect -11089 -388 -11077 388
rect -11043 -388 -11031 388
rect -11089 -400 -11031 -388
rect -10931 388 -10873 400
rect -10931 -388 -10919 388
rect -10885 -388 -10873 388
rect -10931 -400 -10873 -388
rect -10773 388 -10715 400
rect -10773 -388 -10761 388
rect -10727 -388 -10715 388
rect -10773 -400 -10715 -388
rect -10615 388 -10557 400
rect -10615 -388 -10603 388
rect -10569 -388 -10557 388
rect -10615 -400 -10557 -388
rect -10457 388 -10399 400
rect -10457 -388 -10445 388
rect -10411 -388 -10399 388
rect -10457 -400 -10399 -388
rect -10299 388 -10241 400
rect -10299 -388 -10287 388
rect -10253 -388 -10241 388
rect -10299 -400 -10241 -388
rect -10141 388 -10083 400
rect -10141 -388 -10129 388
rect -10095 -388 -10083 388
rect -10141 -400 -10083 -388
rect -9983 388 -9925 400
rect -9983 -388 -9971 388
rect -9937 -388 -9925 388
rect -9983 -400 -9925 -388
rect -9825 388 -9767 400
rect -9825 -388 -9813 388
rect -9779 -388 -9767 388
rect -9825 -400 -9767 -388
rect -9667 388 -9609 400
rect -9667 -388 -9655 388
rect -9621 -388 -9609 388
rect -9667 -400 -9609 -388
rect -9509 388 -9451 400
rect -9509 -388 -9497 388
rect -9463 -388 -9451 388
rect -9509 -400 -9451 -388
rect -9351 388 -9293 400
rect -9351 -388 -9339 388
rect -9305 -388 -9293 388
rect -9351 -400 -9293 -388
rect -9193 388 -9135 400
rect -9193 -388 -9181 388
rect -9147 -388 -9135 388
rect -9193 -400 -9135 -388
rect -9035 388 -8977 400
rect -9035 -388 -9023 388
rect -8989 -388 -8977 388
rect -9035 -400 -8977 -388
rect -8877 388 -8819 400
rect -8877 -388 -8865 388
rect -8831 -388 -8819 388
rect -8877 -400 -8819 -388
rect -8719 388 -8661 400
rect -8719 -388 -8707 388
rect -8673 -388 -8661 388
rect -8719 -400 -8661 -388
rect -8561 388 -8503 400
rect -8561 -388 -8549 388
rect -8515 -388 -8503 388
rect -8561 -400 -8503 -388
rect -8403 388 -8345 400
rect -8403 -388 -8391 388
rect -8357 -388 -8345 388
rect -8403 -400 -8345 -388
rect -8245 388 -8187 400
rect -8245 -388 -8233 388
rect -8199 -388 -8187 388
rect -8245 -400 -8187 -388
rect -8087 388 -8029 400
rect -8087 -388 -8075 388
rect -8041 -388 -8029 388
rect -8087 -400 -8029 -388
rect -7929 388 -7871 400
rect -7929 -388 -7917 388
rect -7883 -388 -7871 388
rect -7929 -400 -7871 -388
rect -7771 388 -7713 400
rect -7771 -388 -7759 388
rect -7725 -388 -7713 388
rect -7771 -400 -7713 -388
rect -7613 388 -7555 400
rect -7613 -388 -7601 388
rect -7567 -388 -7555 388
rect -7613 -400 -7555 -388
rect -7455 388 -7397 400
rect -7455 -388 -7443 388
rect -7409 -388 -7397 388
rect -7455 -400 -7397 -388
rect -7297 388 -7239 400
rect -7297 -388 -7285 388
rect -7251 -388 -7239 388
rect -7297 -400 -7239 -388
rect -7139 388 -7081 400
rect -7139 -388 -7127 388
rect -7093 -388 -7081 388
rect -7139 -400 -7081 -388
rect -6981 388 -6923 400
rect -6981 -388 -6969 388
rect -6935 -388 -6923 388
rect -6981 -400 -6923 -388
rect -6823 388 -6765 400
rect -6823 -388 -6811 388
rect -6777 -388 -6765 388
rect -6823 -400 -6765 -388
rect -6665 388 -6607 400
rect -6665 -388 -6653 388
rect -6619 -388 -6607 388
rect -6665 -400 -6607 -388
rect -6507 388 -6449 400
rect -6507 -388 -6495 388
rect -6461 -388 -6449 388
rect -6507 -400 -6449 -388
rect -6349 388 -6291 400
rect -6349 -388 -6337 388
rect -6303 -388 -6291 388
rect -6349 -400 -6291 -388
rect -6191 388 -6133 400
rect -6191 -388 -6179 388
rect -6145 -388 -6133 388
rect -6191 -400 -6133 -388
rect -6033 388 -5975 400
rect -6033 -388 -6021 388
rect -5987 -388 -5975 388
rect -6033 -400 -5975 -388
rect -5875 388 -5817 400
rect -5875 -388 -5863 388
rect -5829 -388 -5817 388
rect -5875 -400 -5817 -388
rect -5717 388 -5659 400
rect -5717 -388 -5705 388
rect -5671 -388 -5659 388
rect -5717 -400 -5659 -388
rect -5559 388 -5501 400
rect -5559 -388 -5547 388
rect -5513 -388 -5501 388
rect -5559 -400 -5501 -388
rect -5401 388 -5343 400
rect -5401 -388 -5389 388
rect -5355 -388 -5343 388
rect -5401 -400 -5343 -388
rect -5243 388 -5185 400
rect -5243 -388 -5231 388
rect -5197 -388 -5185 388
rect -5243 -400 -5185 -388
rect -5085 388 -5027 400
rect -5085 -388 -5073 388
rect -5039 -388 -5027 388
rect -5085 -400 -5027 -388
rect -4927 388 -4869 400
rect -4927 -388 -4915 388
rect -4881 -388 -4869 388
rect -4927 -400 -4869 -388
rect -4769 388 -4711 400
rect -4769 -388 -4757 388
rect -4723 -388 -4711 388
rect -4769 -400 -4711 -388
rect -4611 388 -4553 400
rect -4611 -388 -4599 388
rect -4565 -388 -4553 388
rect -4611 -400 -4553 -388
rect -4453 388 -4395 400
rect -4453 -388 -4441 388
rect -4407 -388 -4395 388
rect -4453 -400 -4395 -388
rect -4295 388 -4237 400
rect -4295 -388 -4283 388
rect -4249 -388 -4237 388
rect -4295 -400 -4237 -388
rect -4137 388 -4079 400
rect -4137 -388 -4125 388
rect -4091 -388 -4079 388
rect -4137 -400 -4079 -388
rect -3979 388 -3921 400
rect -3979 -388 -3967 388
rect -3933 -388 -3921 388
rect -3979 -400 -3921 -388
rect -3821 388 -3763 400
rect -3821 -388 -3809 388
rect -3775 -388 -3763 388
rect -3821 -400 -3763 -388
rect -3663 388 -3605 400
rect -3663 -388 -3651 388
rect -3617 -388 -3605 388
rect -3663 -400 -3605 -388
rect -3505 388 -3447 400
rect -3505 -388 -3493 388
rect -3459 -388 -3447 388
rect -3505 -400 -3447 -388
rect -3347 388 -3289 400
rect -3347 -388 -3335 388
rect -3301 -388 -3289 388
rect -3347 -400 -3289 -388
rect -3189 388 -3131 400
rect -3189 -388 -3177 388
rect -3143 -388 -3131 388
rect -3189 -400 -3131 -388
rect -3031 388 -2973 400
rect -3031 -388 -3019 388
rect -2985 -388 -2973 388
rect -3031 -400 -2973 -388
rect -2873 388 -2815 400
rect -2873 -388 -2861 388
rect -2827 -388 -2815 388
rect -2873 -400 -2815 -388
rect -2715 388 -2657 400
rect -2715 -388 -2703 388
rect -2669 -388 -2657 388
rect -2715 -400 -2657 -388
rect -2557 388 -2499 400
rect -2557 -388 -2545 388
rect -2511 -388 -2499 388
rect -2557 -400 -2499 -388
rect -2399 388 -2341 400
rect -2399 -388 -2387 388
rect -2353 -388 -2341 388
rect -2399 -400 -2341 -388
rect -2241 388 -2183 400
rect -2241 -388 -2229 388
rect -2195 -388 -2183 388
rect -2241 -400 -2183 -388
rect -2083 388 -2025 400
rect -2083 -388 -2071 388
rect -2037 -388 -2025 388
rect -2083 -400 -2025 -388
rect -1925 388 -1867 400
rect -1925 -388 -1913 388
rect -1879 -388 -1867 388
rect -1925 -400 -1867 -388
rect -1767 388 -1709 400
rect -1767 -388 -1755 388
rect -1721 -388 -1709 388
rect -1767 -400 -1709 -388
rect -1609 388 -1551 400
rect -1609 -388 -1597 388
rect -1563 -388 -1551 388
rect -1609 -400 -1551 -388
rect -1451 388 -1393 400
rect -1451 -388 -1439 388
rect -1405 -388 -1393 388
rect -1451 -400 -1393 -388
rect -1293 388 -1235 400
rect -1293 -388 -1281 388
rect -1247 -388 -1235 388
rect -1293 -400 -1235 -388
rect -1135 388 -1077 400
rect -1135 -388 -1123 388
rect -1089 -388 -1077 388
rect -1135 -400 -1077 -388
rect -977 388 -919 400
rect -977 -388 -965 388
rect -931 -388 -919 388
rect -977 -400 -919 -388
rect -819 388 -761 400
rect -819 -388 -807 388
rect -773 -388 -761 388
rect -819 -400 -761 -388
rect -661 388 -603 400
rect -661 -388 -649 388
rect -615 -388 -603 388
rect -661 -400 -603 -388
rect -503 388 -445 400
rect -503 -388 -491 388
rect -457 -388 -445 388
rect -503 -400 -445 -388
rect -345 388 -287 400
rect -345 -388 -333 388
rect -299 -388 -287 388
rect -345 -400 -287 -388
rect -187 388 -129 400
rect -187 -388 -175 388
rect -141 -388 -129 388
rect -187 -400 -129 -388
rect -29 388 29 400
rect -29 -388 -17 388
rect 17 -388 29 388
rect -29 -400 29 -388
rect 129 388 187 400
rect 129 -388 141 388
rect 175 -388 187 388
rect 129 -400 187 -388
rect 287 388 345 400
rect 287 -388 299 388
rect 333 -388 345 388
rect 287 -400 345 -388
rect 445 388 503 400
rect 445 -388 457 388
rect 491 -388 503 388
rect 445 -400 503 -388
rect 603 388 661 400
rect 603 -388 615 388
rect 649 -388 661 388
rect 603 -400 661 -388
rect 761 388 819 400
rect 761 -388 773 388
rect 807 -388 819 388
rect 761 -400 819 -388
rect 919 388 977 400
rect 919 -388 931 388
rect 965 -388 977 388
rect 919 -400 977 -388
rect 1077 388 1135 400
rect 1077 -388 1089 388
rect 1123 -388 1135 388
rect 1077 -400 1135 -388
rect 1235 388 1293 400
rect 1235 -388 1247 388
rect 1281 -388 1293 388
rect 1235 -400 1293 -388
rect 1393 388 1451 400
rect 1393 -388 1405 388
rect 1439 -388 1451 388
rect 1393 -400 1451 -388
rect 1551 388 1609 400
rect 1551 -388 1563 388
rect 1597 -388 1609 388
rect 1551 -400 1609 -388
rect 1709 388 1767 400
rect 1709 -388 1721 388
rect 1755 -388 1767 388
rect 1709 -400 1767 -388
rect 1867 388 1925 400
rect 1867 -388 1879 388
rect 1913 -388 1925 388
rect 1867 -400 1925 -388
rect 2025 388 2083 400
rect 2025 -388 2037 388
rect 2071 -388 2083 388
rect 2025 -400 2083 -388
rect 2183 388 2241 400
rect 2183 -388 2195 388
rect 2229 -388 2241 388
rect 2183 -400 2241 -388
rect 2341 388 2399 400
rect 2341 -388 2353 388
rect 2387 -388 2399 388
rect 2341 -400 2399 -388
rect 2499 388 2557 400
rect 2499 -388 2511 388
rect 2545 -388 2557 388
rect 2499 -400 2557 -388
rect 2657 388 2715 400
rect 2657 -388 2669 388
rect 2703 -388 2715 388
rect 2657 -400 2715 -388
rect 2815 388 2873 400
rect 2815 -388 2827 388
rect 2861 -388 2873 388
rect 2815 -400 2873 -388
rect 2973 388 3031 400
rect 2973 -388 2985 388
rect 3019 -388 3031 388
rect 2973 -400 3031 -388
rect 3131 388 3189 400
rect 3131 -388 3143 388
rect 3177 -388 3189 388
rect 3131 -400 3189 -388
rect 3289 388 3347 400
rect 3289 -388 3301 388
rect 3335 -388 3347 388
rect 3289 -400 3347 -388
rect 3447 388 3505 400
rect 3447 -388 3459 388
rect 3493 -388 3505 388
rect 3447 -400 3505 -388
rect 3605 388 3663 400
rect 3605 -388 3617 388
rect 3651 -388 3663 388
rect 3605 -400 3663 -388
rect 3763 388 3821 400
rect 3763 -388 3775 388
rect 3809 -388 3821 388
rect 3763 -400 3821 -388
rect 3921 388 3979 400
rect 3921 -388 3933 388
rect 3967 -388 3979 388
rect 3921 -400 3979 -388
rect 4079 388 4137 400
rect 4079 -388 4091 388
rect 4125 -388 4137 388
rect 4079 -400 4137 -388
rect 4237 388 4295 400
rect 4237 -388 4249 388
rect 4283 -388 4295 388
rect 4237 -400 4295 -388
rect 4395 388 4453 400
rect 4395 -388 4407 388
rect 4441 -388 4453 388
rect 4395 -400 4453 -388
rect 4553 388 4611 400
rect 4553 -388 4565 388
rect 4599 -388 4611 388
rect 4553 -400 4611 -388
rect 4711 388 4769 400
rect 4711 -388 4723 388
rect 4757 -388 4769 388
rect 4711 -400 4769 -388
rect 4869 388 4927 400
rect 4869 -388 4881 388
rect 4915 -388 4927 388
rect 4869 -400 4927 -388
rect 5027 388 5085 400
rect 5027 -388 5039 388
rect 5073 -388 5085 388
rect 5027 -400 5085 -388
rect 5185 388 5243 400
rect 5185 -388 5197 388
rect 5231 -388 5243 388
rect 5185 -400 5243 -388
rect 5343 388 5401 400
rect 5343 -388 5355 388
rect 5389 -388 5401 388
rect 5343 -400 5401 -388
rect 5501 388 5559 400
rect 5501 -388 5513 388
rect 5547 -388 5559 388
rect 5501 -400 5559 -388
rect 5659 388 5717 400
rect 5659 -388 5671 388
rect 5705 -388 5717 388
rect 5659 -400 5717 -388
rect 5817 388 5875 400
rect 5817 -388 5829 388
rect 5863 -388 5875 388
rect 5817 -400 5875 -388
rect 5975 388 6033 400
rect 5975 -388 5987 388
rect 6021 -388 6033 388
rect 5975 -400 6033 -388
rect 6133 388 6191 400
rect 6133 -388 6145 388
rect 6179 -388 6191 388
rect 6133 -400 6191 -388
rect 6291 388 6349 400
rect 6291 -388 6303 388
rect 6337 -388 6349 388
rect 6291 -400 6349 -388
rect 6449 388 6507 400
rect 6449 -388 6461 388
rect 6495 -388 6507 388
rect 6449 -400 6507 -388
rect 6607 388 6665 400
rect 6607 -388 6619 388
rect 6653 -388 6665 388
rect 6607 -400 6665 -388
rect 6765 388 6823 400
rect 6765 -388 6777 388
rect 6811 -388 6823 388
rect 6765 -400 6823 -388
rect 6923 388 6981 400
rect 6923 -388 6935 388
rect 6969 -388 6981 388
rect 6923 -400 6981 -388
rect 7081 388 7139 400
rect 7081 -388 7093 388
rect 7127 -388 7139 388
rect 7081 -400 7139 -388
rect 7239 388 7297 400
rect 7239 -388 7251 388
rect 7285 -388 7297 388
rect 7239 -400 7297 -388
rect 7397 388 7455 400
rect 7397 -388 7409 388
rect 7443 -388 7455 388
rect 7397 -400 7455 -388
rect 7555 388 7613 400
rect 7555 -388 7567 388
rect 7601 -388 7613 388
rect 7555 -400 7613 -388
rect 7713 388 7771 400
rect 7713 -388 7725 388
rect 7759 -388 7771 388
rect 7713 -400 7771 -388
rect 7871 388 7929 400
rect 7871 -388 7883 388
rect 7917 -388 7929 388
rect 7871 -400 7929 -388
rect 8029 388 8087 400
rect 8029 -388 8041 388
rect 8075 -388 8087 388
rect 8029 -400 8087 -388
rect 8187 388 8245 400
rect 8187 -388 8199 388
rect 8233 -388 8245 388
rect 8187 -400 8245 -388
rect 8345 388 8403 400
rect 8345 -388 8357 388
rect 8391 -388 8403 388
rect 8345 -400 8403 -388
rect 8503 388 8561 400
rect 8503 -388 8515 388
rect 8549 -388 8561 388
rect 8503 -400 8561 -388
rect 8661 388 8719 400
rect 8661 -388 8673 388
rect 8707 -388 8719 388
rect 8661 -400 8719 -388
rect 8819 388 8877 400
rect 8819 -388 8831 388
rect 8865 -388 8877 388
rect 8819 -400 8877 -388
rect 8977 388 9035 400
rect 8977 -388 8989 388
rect 9023 -388 9035 388
rect 8977 -400 9035 -388
rect 9135 388 9193 400
rect 9135 -388 9147 388
rect 9181 -388 9193 388
rect 9135 -400 9193 -388
rect 9293 388 9351 400
rect 9293 -388 9305 388
rect 9339 -388 9351 388
rect 9293 -400 9351 -388
rect 9451 388 9509 400
rect 9451 -388 9463 388
rect 9497 -388 9509 388
rect 9451 -400 9509 -388
rect 9609 388 9667 400
rect 9609 -388 9621 388
rect 9655 -388 9667 388
rect 9609 -400 9667 -388
rect 9767 388 9825 400
rect 9767 -388 9779 388
rect 9813 -388 9825 388
rect 9767 -400 9825 -388
rect 9925 388 9983 400
rect 9925 -388 9937 388
rect 9971 -388 9983 388
rect 9925 -400 9983 -388
rect 10083 388 10141 400
rect 10083 -388 10095 388
rect 10129 -388 10141 388
rect 10083 -400 10141 -388
rect 10241 388 10299 400
rect 10241 -388 10253 388
rect 10287 -388 10299 388
rect 10241 -400 10299 -388
rect 10399 388 10457 400
rect 10399 -388 10411 388
rect 10445 -388 10457 388
rect 10399 -400 10457 -388
rect 10557 388 10615 400
rect 10557 -388 10569 388
rect 10603 -388 10615 388
rect 10557 -400 10615 -388
rect 10715 388 10773 400
rect 10715 -388 10727 388
rect 10761 -388 10773 388
rect 10715 -400 10773 -388
rect 10873 388 10931 400
rect 10873 -388 10885 388
rect 10919 -388 10931 388
rect 10873 -400 10931 -388
rect 11031 388 11089 400
rect 11031 -388 11043 388
rect 11077 -388 11089 388
rect 11031 -400 11089 -388
rect 11189 388 11247 400
rect 11189 -388 11201 388
rect 11235 -388 11247 388
rect 11189 -400 11247 -388
rect 11347 388 11405 400
rect 11347 -388 11359 388
rect 11393 -388 11405 388
rect 11347 -400 11405 -388
rect 11505 388 11563 400
rect 11505 -388 11517 388
rect 11551 -388 11563 388
rect 11505 -400 11563 -388
rect 11663 388 11721 400
rect 11663 -388 11675 388
rect 11709 -388 11721 388
rect 11663 -400 11721 -388
rect 11821 388 11879 400
rect 11821 -388 11833 388
rect 11867 -388 11879 388
rect 11821 -400 11879 -388
rect 11979 388 12037 400
rect 11979 -388 11991 388
rect 12025 -388 12037 388
rect 11979 -400 12037 -388
rect 12137 388 12195 400
rect 12137 -388 12149 388
rect 12183 -388 12195 388
rect 12137 -400 12195 -388
rect 12295 388 12353 400
rect 12295 -388 12307 388
rect 12341 -388 12353 388
rect 12295 -400 12353 -388
rect 12453 388 12511 400
rect 12453 -388 12465 388
rect 12499 -388 12511 388
rect 12453 -400 12511 -388
rect 12611 388 12669 400
rect 12611 -388 12623 388
rect 12657 -388 12669 388
rect 12611 -400 12669 -388
rect 12769 388 12827 400
rect 12769 -388 12781 388
rect 12815 -388 12827 388
rect 12769 -400 12827 -388
rect 12927 388 12985 400
rect 12927 -388 12939 388
rect 12973 -388 12985 388
rect 12927 -400 12985 -388
<< mvndiffc >>
rect -12973 -388 -12939 388
rect -12815 -388 -12781 388
rect -12657 -388 -12623 388
rect -12499 -388 -12465 388
rect -12341 -388 -12307 388
rect -12183 -388 -12149 388
rect -12025 -388 -11991 388
rect -11867 -388 -11833 388
rect -11709 -388 -11675 388
rect -11551 -388 -11517 388
rect -11393 -388 -11359 388
rect -11235 -388 -11201 388
rect -11077 -388 -11043 388
rect -10919 -388 -10885 388
rect -10761 -388 -10727 388
rect -10603 -388 -10569 388
rect -10445 -388 -10411 388
rect -10287 -388 -10253 388
rect -10129 -388 -10095 388
rect -9971 -388 -9937 388
rect -9813 -388 -9779 388
rect -9655 -388 -9621 388
rect -9497 -388 -9463 388
rect -9339 -388 -9305 388
rect -9181 -388 -9147 388
rect -9023 -388 -8989 388
rect -8865 -388 -8831 388
rect -8707 -388 -8673 388
rect -8549 -388 -8515 388
rect -8391 -388 -8357 388
rect -8233 -388 -8199 388
rect -8075 -388 -8041 388
rect -7917 -388 -7883 388
rect -7759 -388 -7725 388
rect -7601 -388 -7567 388
rect -7443 -388 -7409 388
rect -7285 -388 -7251 388
rect -7127 -388 -7093 388
rect -6969 -388 -6935 388
rect -6811 -388 -6777 388
rect -6653 -388 -6619 388
rect -6495 -388 -6461 388
rect -6337 -388 -6303 388
rect -6179 -388 -6145 388
rect -6021 -388 -5987 388
rect -5863 -388 -5829 388
rect -5705 -388 -5671 388
rect -5547 -388 -5513 388
rect -5389 -388 -5355 388
rect -5231 -388 -5197 388
rect -5073 -388 -5039 388
rect -4915 -388 -4881 388
rect -4757 -388 -4723 388
rect -4599 -388 -4565 388
rect -4441 -388 -4407 388
rect -4283 -388 -4249 388
rect -4125 -388 -4091 388
rect -3967 -388 -3933 388
rect -3809 -388 -3775 388
rect -3651 -388 -3617 388
rect -3493 -388 -3459 388
rect -3335 -388 -3301 388
rect -3177 -388 -3143 388
rect -3019 -388 -2985 388
rect -2861 -388 -2827 388
rect -2703 -388 -2669 388
rect -2545 -388 -2511 388
rect -2387 -388 -2353 388
rect -2229 -388 -2195 388
rect -2071 -388 -2037 388
rect -1913 -388 -1879 388
rect -1755 -388 -1721 388
rect -1597 -388 -1563 388
rect -1439 -388 -1405 388
rect -1281 -388 -1247 388
rect -1123 -388 -1089 388
rect -965 -388 -931 388
rect -807 -388 -773 388
rect -649 -388 -615 388
rect -491 -388 -457 388
rect -333 -388 -299 388
rect -175 -388 -141 388
rect -17 -388 17 388
rect 141 -388 175 388
rect 299 -388 333 388
rect 457 -388 491 388
rect 615 -388 649 388
rect 773 -388 807 388
rect 931 -388 965 388
rect 1089 -388 1123 388
rect 1247 -388 1281 388
rect 1405 -388 1439 388
rect 1563 -388 1597 388
rect 1721 -388 1755 388
rect 1879 -388 1913 388
rect 2037 -388 2071 388
rect 2195 -388 2229 388
rect 2353 -388 2387 388
rect 2511 -388 2545 388
rect 2669 -388 2703 388
rect 2827 -388 2861 388
rect 2985 -388 3019 388
rect 3143 -388 3177 388
rect 3301 -388 3335 388
rect 3459 -388 3493 388
rect 3617 -388 3651 388
rect 3775 -388 3809 388
rect 3933 -388 3967 388
rect 4091 -388 4125 388
rect 4249 -388 4283 388
rect 4407 -388 4441 388
rect 4565 -388 4599 388
rect 4723 -388 4757 388
rect 4881 -388 4915 388
rect 5039 -388 5073 388
rect 5197 -388 5231 388
rect 5355 -388 5389 388
rect 5513 -388 5547 388
rect 5671 -388 5705 388
rect 5829 -388 5863 388
rect 5987 -388 6021 388
rect 6145 -388 6179 388
rect 6303 -388 6337 388
rect 6461 -388 6495 388
rect 6619 -388 6653 388
rect 6777 -388 6811 388
rect 6935 -388 6969 388
rect 7093 -388 7127 388
rect 7251 -388 7285 388
rect 7409 -388 7443 388
rect 7567 -388 7601 388
rect 7725 -388 7759 388
rect 7883 -388 7917 388
rect 8041 -388 8075 388
rect 8199 -388 8233 388
rect 8357 -388 8391 388
rect 8515 -388 8549 388
rect 8673 -388 8707 388
rect 8831 -388 8865 388
rect 8989 -388 9023 388
rect 9147 -388 9181 388
rect 9305 -388 9339 388
rect 9463 -388 9497 388
rect 9621 -388 9655 388
rect 9779 -388 9813 388
rect 9937 -388 9971 388
rect 10095 -388 10129 388
rect 10253 -388 10287 388
rect 10411 -388 10445 388
rect 10569 -388 10603 388
rect 10727 -388 10761 388
rect 10885 -388 10919 388
rect 11043 -388 11077 388
rect 11201 -388 11235 388
rect 11359 -388 11393 388
rect 11517 -388 11551 388
rect 11675 -388 11709 388
rect 11833 -388 11867 388
rect 11991 -388 12025 388
rect 12149 -388 12183 388
rect 12307 -388 12341 388
rect 12465 -388 12499 388
rect 12623 -388 12657 388
rect 12781 -388 12815 388
rect 12939 -388 12973 388
<< mvpsubdiff >>
rect -13119 610 13119 622
rect -13119 576 -13011 610
rect 13011 576 13119 610
rect -13119 564 13119 576
rect -13119 514 -13061 564
rect -13119 -514 -13107 514
rect -13073 -514 -13061 514
rect 13061 514 13119 564
rect -13119 -564 -13061 -514
rect 13061 -514 13073 514
rect 13107 -514 13119 514
rect 13061 -564 13119 -514
rect -13119 -576 13119 -564
rect -13119 -610 -13011 -576
rect 13011 -610 13119 -576
rect -13119 -622 13119 -610
<< mvpsubdiffcont >>
rect -13011 576 13011 610
rect -13107 -514 -13073 514
rect 13073 -514 13107 514
rect -13011 -610 13011 -576
<< poly >>
rect -12927 472 -12827 488
rect -12927 438 -12911 472
rect -12843 438 -12827 472
rect -12927 400 -12827 438
rect -12769 472 -12669 488
rect -12769 438 -12753 472
rect -12685 438 -12669 472
rect -12769 400 -12669 438
rect -12611 472 -12511 488
rect -12611 438 -12595 472
rect -12527 438 -12511 472
rect -12611 400 -12511 438
rect -12453 472 -12353 488
rect -12453 438 -12437 472
rect -12369 438 -12353 472
rect -12453 400 -12353 438
rect -12295 472 -12195 488
rect -12295 438 -12279 472
rect -12211 438 -12195 472
rect -12295 400 -12195 438
rect -12137 472 -12037 488
rect -12137 438 -12121 472
rect -12053 438 -12037 472
rect -12137 400 -12037 438
rect -11979 472 -11879 488
rect -11979 438 -11963 472
rect -11895 438 -11879 472
rect -11979 400 -11879 438
rect -11821 472 -11721 488
rect -11821 438 -11805 472
rect -11737 438 -11721 472
rect -11821 400 -11721 438
rect -11663 472 -11563 488
rect -11663 438 -11647 472
rect -11579 438 -11563 472
rect -11663 400 -11563 438
rect -11505 472 -11405 488
rect -11505 438 -11489 472
rect -11421 438 -11405 472
rect -11505 400 -11405 438
rect -11347 472 -11247 488
rect -11347 438 -11331 472
rect -11263 438 -11247 472
rect -11347 400 -11247 438
rect -11189 472 -11089 488
rect -11189 438 -11173 472
rect -11105 438 -11089 472
rect -11189 400 -11089 438
rect -11031 472 -10931 488
rect -11031 438 -11015 472
rect -10947 438 -10931 472
rect -11031 400 -10931 438
rect -10873 472 -10773 488
rect -10873 438 -10857 472
rect -10789 438 -10773 472
rect -10873 400 -10773 438
rect -10715 472 -10615 488
rect -10715 438 -10699 472
rect -10631 438 -10615 472
rect -10715 400 -10615 438
rect -10557 472 -10457 488
rect -10557 438 -10541 472
rect -10473 438 -10457 472
rect -10557 400 -10457 438
rect -10399 472 -10299 488
rect -10399 438 -10383 472
rect -10315 438 -10299 472
rect -10399 400 -10299 438
rect -10241 472 -10141 488
rect -10241 438 -10225 472
rect -10157 438 -10141 472
rect -10241 400 -10141 438
rect -10083 472 -9983 488
rect -10083 438 -10067 472
rect -9999 438 -9983 472
rect -10083 400 -9983 438
rect -9925 472 -9825 488
rect -9925 438 -9909 472
rect -9841 438 -9825 472
rect -9925 400 -9825 438
rect -9767 472 -9667 488
rect -9767 438 -9751 472
rect -9683 438 -9667 472
rect -9767 400 -9667 438
rect -9609 472 -9509 488
rect -9609 438 -9593 472
rect -9525 438 -9509 472
rect -9609 400 -9509 438
rect -9451 472 -9351 488
rect -9451 438 -9435 472
rect -9367 438 -9351 472
rect -9451 400 -9351 438
rect -9293 472 -9193 488
rect -9293 438 -9277 472
rect -9209 438 -9193 472
rect -9293 400 -9193 438
rect -9135 472 -9035 488
rect -9135 438 -9119 472
rect -9051 438 -9035 472
rect -9135 400 -9035 438
rect -8977 472 -8877 488
rect -8977 438 -8961 472
rect -8893 438 -8877 472
rect -8977 400 -8877 438
rect -8819 472 -8719 488
rect -8819 438 -8803 472
rect -8735 438 -8719 472
rect -8819 400 -8719 438
rect -8661 472 -8561 488
rect -8661 438 -8645 472
rect -8577 438 -8561 472
rect -8661 400 -8561 438
rect -8503 472 -8403 488
rect -8503 438 -8487 472
rect -8419 438 -8403 472
rect -8503 400 -8403 438
rect -8345 472 -8245 488
rect -8345 438 -8329 472
rect -8261 438 -8245 472
rect -8345 400 -8245 438
rect -8187 472 -8087 488
rect -8187 438 -8171 472
rect -8103 438 -8087 472
rect -8187 400 -8087 438
rect -8029 472 -7929 488
rect -8029 438 -8013 472
rect -7945 438 -7929 472
rect -8029 400 -7929 438
rect -7871 472 -7771 488
rect -7871 438 -7855 472
rect -7787 438 -7771 472
rect -7871 400 -7771 438
rect -7713 472 -7613 488
rect -7713 438 -7697 472
rect -7629 438 -7613 472
rect -7713 400 -7613 438
rect -7555 472 -7455 488
rect -7555 438 -7539 472
rect -7471 438 -7455 472
rect -7555 400 -7455 438
rect -7397 472 -7297 488
rect -7397 438 -7381 472
rect -7313 438 -7297 472
rect -7397 400 -7297 438
rect -7239 472 -7139 488
rect -7239 438 -7223 472
rect -7155 438 -7139 472
rect -7239 400 -7139 438
rect -7081 472 -6981 488
rect -7081 438 -7065 472
rect -6997 438 -6981 472
rect -7081 400 -6981 438
rect -6923 472 -6823 488
rect -6923 438 -6907 472
rect -6839 438 -6823 472
rect -6923 400 -6823 438
rect -6765 472 -6665 488
rect -6765 438 -6749 472
rect -6681 438 -6665 472
rect -6765 400 -6665 438
rect -6607 472 -6507 488
rect -6607 438 -6591 472
rect -6523 438 -6507 472
rect -6607 400 -6507 438
rect -6449 472 -6349 488
rect -6449 438 -6433 472
rect -6365 438 -6349 472
rect -6449 400 -6349 438
rect -6291 472 -6191 488
rect -6291 438 -6275 472
rect -6207 438 -6191 472
rect -6291 400 -6191 438
rect -6133 472 -6033 488
rect -6133 438 -6117 472
rect -6049 438 -6033 472
rect -6133 400 -6033 438
rect -5975 472 -5875 488
rect -5975 438 -5959 472
rect -5891 438 -5875 472
rect -5975 400 -5875 438
rect -5817 472 -5717 488
rect -5817 438 -5801 472
rect -5733 438 -5717 472
rect -5817 400 -5717 438
rect -5659 472 -5559 488
rect -5659 438 -5643 472
rect -5575 438 -5559 472
rect -5659 400 -5559 438
rect -5501 472 -5401 488
rect -5501 438 -5485 472
rect -5417 438 -5401 472
rect -5501 400 -5401 438
rect -5343 472 -5243 488
rect -5343 438 -5327 472
rect -5259 438 -5243 472
rect -5343 400 -5243 438
rect -5185 472 -5085 488
rect -5185 438 -5169 472
rect -5101 438 -5085 472
rect -5185 400 -5085 438
rect -5027 472 -4927 488
rect -5027 438 -5011 472
rect -4943 438 -4927 472
rect -5027 400 -4927 438
rect -4869 472 -4769 488
rect -4869 438 -4853 472
rect -4785 438 -4769 472
rect -4869 400 -4769 438
rect -4711 472 -4611 488
rect -4711 438 -4695 472
rect -4627 438 -4611 472
rect -4711 400 -4611 438
rect -4553 472 -4453 488
rect -4553 438 -4537 472
rect -4469 438 -4453 472
rect -4553 400 -4453 438
rect -4395 472 -4295 488
rect -4395 438 -4379 472
rect -4311 438 -4295 472
rect -4395 400 -4295 438
rect -4237 472 -4137 488
rect -4237 438 -4221 472
rect -4153 438 -4137 472
rect -4237 400 -4137 438
rect -4079 472 -3979 488
rect -4079 438 -4063 472
rect -3995 438 -3979 472
rect -4079 400 -3979 438
rect -3921 472 -3821 488
rect -3921 438 -3905 472
rect -3837 438 -3821 472
rect -3921 400 -3821 438
rect -3763 472 -3663 488
rect -3763 438 -3747 472
rect -3679 438 -3663 472
rect -3763 400 -3663 438
rect -3605 472 -3505 488
rect -3605 438 -3589 472
rect -3521 438 -3505 472
rect -3605 400 -3505 438
rect -3447 472 -3347 488
rect -3447 438 -3431 472
rect -3363 438 -3347 472
rect -3447 400 -3347 438
rect -3289 472 -3189 488
rect -3289 438 -3273 472
rect -3205 438 -3189 472
rect -3289 400 -3189 438
rect -3131 472 -3031 488
rect -3131 438 -3115 472
rect -3047 438 -3031 472
rect -3131 400 -3031 438
rect -2973 472 -2873 488
rect -2973 438 -2957 472
rect -2889 438 -2873 472
rect -2973 400 -2873 438
rect -2815 472 -2715 488
rect -2815 438 -2799 472
rect -2731 438 -2715 472
rect -2815 400 -2715 438
rect -2657 472 -2557 488
rect -2657 438 -2641 472
rect -2573 438 -2557 472
rect -2657 400 -2557 438
rect -2499 472 -2399 488
rect -2499 438 -2483 472
rect -2415 438 -2399 472
rect -2499 400 -2399 438
rect -2341 472 -2241 488
rect -2341 438 -2325 472
rect -2257 438 -2241 472
rect -2341 400 -2241 438
rect -2183 472 -2083 488
rect -2183 438 -2167 472
rect -2099 438 -2083 472
rect -2183 400 -2083 438
rect -2025 472 -1925 488
rect -2025 438 -2009 472
rect -1941 438 -1925 472
rect -2025 400 -1925 438
rect -1867 472 -1767 488
rect -1867 438 -1851 472
rect -1783 438 -1767 472
rect -1867 400 -1767 438
rect -1709 472 -1609 488
rect -1709 438 -1693 472
rect -1625 438 -1609 472
rect -1709 400 -1609 438
rect -1551 472 -1451 488
rect -1551 438 -1535 472
rect -1467 438 -1451 472
rect -1551 400 -1451 438
rect -1393 472 -1293 488
rect -1393 438 -1377 472
rect -1309 438 -1293 472
rect -1393 400 -1293 438
rect -1235 472 -1135 488
rect -1235 438 -1219 472
rect -1151 438 -1135 472
rect -1235 400 -1135 438
rect -1077 472 -977 488
rect -1077 438 -1061 472
rect -993 438 -977 472
rect -1077 400 -977 438
rect -919 472 -819 488
rect -919 438 -903 472
rect -835 438 -819 472
rect -919 400 -819 438
rect -761 472 -661 488
rect -761 438 -745 472
rect -677 438 -661 472
rect -761 400 -661 438
rect -603 472 -503 488
rect -603 438 -587 472
rect -519 438 -503 472
rect -603 400 -503 438
rect -445 472 -345 488
rect -445 438 -429 472
rect -361 438 -345 472
rect -445 400 -345 438
rect -287 472 -187 488
rect -287 438 -271 472
rect -203 438 -187 472
rect -287 400 -187 438
rect -129 472 -29 488
rect -129 438 -113 472
rect -45 438 -29 472
rect -129 400 -29 438
rect 29 472 129 488
rect 29 438 45 472
rect 113 438 129 472
rect 29 400 129 438
rect 187 472 287 488
rect 187 438 203 472
rect 271 438 287 472
rect 187 400 287 438
rect 345 472 445 488
rect 345 438 361 472
rect 429 438 445 472
rect 345 400 445 438
rect 503 472 603 488
rect 503 438 519 472
rect 587 438 603 472
rect 503 400 603 438
rect 661 472 761 488
rect 661 438 677 472
rect 745 438 761 472
rect 661 400 761 438
rect 819 472 919 488
rect 819 438 835 472
rect 903 438 919 472
rect 819 400 919 438
rect 977 472 1077 488
rect 977 438 993 472
rect 1061 438 1077 472
rect 977 400 1077 438
rect 1135 472 1235 488
rect 1135 438 1151 472
rect 1219 438 1235 472
rect 1135 400 1235 438
rect 1293 472 1393 488
rect 1293 438 1309 472
rect 1377 438 1393 472
rect 1293 400 1393 438
rect 1451 472 1551 488
rect 1451 438 1467 472
rect 1535 438 1551 472
rect 1451 400 1551 438
rect 1609 472 1709 488
rect 1609 438 1625 472
rect 1693 438 1709 472
rect 1609 400 1709 438
rect 1767 472 1867 488
rect 1767 438 1783 472
rect 1851 438 1867 472
rect 1767 400 1867 438
rect 1925 472 2025 488
rect 1925 438 1941 472
rect 2009 438 2025 472
rect 1925 400 2025 438
rect 2083 472 2183 488
rect 2083 438 2099 472
rect 2167 438 2183 472
rect 2083 400 2183 438
rect 2241 472 2341 488
rect 2241 438 2257 472
rect 2325 438 2341 472
rect 2241 400 2341 438
rect 2399 472 2499 488
rect 2399 438 2415 472
rect 2483 438 2499 472
rect 2399 400 2499 438
rect 2557 472 2657 488
rect 2557 438 2573 472
rect 2641 438 2657 472
rect 2557 400 2657 438
rect 2715 472 2815 488
rect 2715 438 2731 472
rect 2799 438 2815 472
rect 2715 400 2815 438
rect 2873 472 2973 488
rect 2873 438 2889 472
rect 2957 438 2973 472
rect 2873 400 2973 438
rect 3031 472 3131 488
rect 3031 438 3047 472
rect 3115 438 3131 472
rect 3031 400 3131 438
rect 3189 472 3289 488
rect 3189 438 3205 472
rect 3273 438 3289 472
rect 3189 400 3289 438
rect 3347 472 3447 488
rect 3347 438 3363 472
rect 3431 438 3447 472
rect 3347 400 3447 438
rect 3505 472 3605 488
rect 3505 438 3521 472
rect 3589 438 3605 472
rect 3505 400 3605 438
rect 3663 472 3763 488
rect 3663 438 3679 472
rect 3747 438 3763 472
rect 3663 400 3763 438
rect 3821 472 3921 488
rect 3821 438 3837 472
rect 3905 438 3921 472
rect 3821 400 3921 438
rect 3979 472 4079 488
rect 3979 438 3995 472
rect 4063 438 4079 472
rect 3979 400 4079 438
rect 4137 472 4237 488
rect 4137 438 4153 472
rect 4221 438 4237 472
rect 4137 400 4237 438
rect 4295 472 4395 488
rect 4295 438 4311 472
rect 4379 438 4395 472
rect 4295 400 4395 438
rect 4453 472 4553 488
rect 4453 438 4469 472
rect 4537 438 4553 472
rect 4453 400 4553 438
rect 4611 472 4711 488
rect 4611 438 4627 472
rect 4695 438 4711 472
rect 4611 400 4711 438
rect 4769 472 4869 488
rect 4769 438 4785 472
rect 4853 438 4869 472
rect 4769 400 4869 438
rect 4927 472 5027 488
rect 4927 438 4943 472
rect 5011 438 5027 472
rect 4927 400 5027 438
rect 5085 472 5185 488
rect 5085 438 5101 472
rect 5169 438 5185 472
rect 5085 400 5185 438
rect 5243 472 5343 488
rect 5243 438 5259 472
rect 5327 438 5343 472
rect 5243 400 5343 438
rect 5401 472 5501 488
rect 5401 438 5417 472
rect 5485 438 5501 472
rect 5401 400 5501 438
rect 5559 472 5659 488
rect 5559 438 5575 472
rect 5643 438 5659 472
rect 5559 400 5659 438
rect 5717 472 5817 488
rect 5717 438 5733 472
rect 5801 438 5817 472
rect 5717 400 5817 438
rect 5875 472 5975 488
rect 5875 438 5891 472
rect 5959 438 5975 472
rect 5875 400 5975 438
rect 6033 472 6133 488
rect 6033 438 6049 472
rect 6117 438 6133 472
rect 6033 400 6133 438
rect 6191 472 6291 488
rect 6191 438 6207 472
rect 6275 438 6291 472
rect 6191 400 6291 438
rect 6349 472 6449 488
rect 6349 438 6365 472
rect 6433 438 6449 472
rect 6349 400 6449 438
rect 6507 472 6607 488
rect 6507 438 6523 472
rect 6591 438 6607 472
rect 6507 400 6607 438
rect 6665 472 6765 488
rect 6665 438 6681 472
rect 6749 438 6765 472
rect 6665 400 6765 438
rect 6823 472 6923 488
rect 6823 438 6839 472
rect 6907 438 6923 472
rect 6823 400 6923 438
rect 6981 472 7081 488
rect 6981 438 6997 472
rect 7065 438 7081 472
rect 6981 400 7081 438
rect 7139 472 7239 488
rect 7139 438 7155 472
rect 7223 438 7239 472
rect 7139 400 7239 438
rect 7297 472 7397 488
rect 7297 438 7313 472
rect 7381 438 7397 472
rect 7297 400 7397 438
rect 7455 472 7555 488
rect 7455 438 7471 472
rect 7539 438 7555 472
rect 7455 400 7555 438
rect 7613 472 7713 488
rect 7613 438 7629 472
rect 7697 438 7713 472
rect 7613 400 7713 438
rect 7771 472 7871 488
rect 7771 438 7787 472
rect 7855 438 7871 472
rect 7771 400 7871 438
rect 7929 472 8029 488
rect 7929 438 7945 472
rect 8013 438 8029 472
rect 7929 400 8029 438
rect 8087 472 8187 488
rect 8087 438 8103 472
rect 8171 438 8187 472
rect 8087 400 8187 438
rect 8245 472 8345 488
rect 8245 438 8261 472
rect 8329 438 8345 472
rect 8245 400 8345 438
rect 8403 472 8503 488
rect 8403 438 8419 472
rect 8487 438 8503 472
rect 8403 400 8503 438
rect 8561 472 8661 488
rect 8561 438 8577 472
rect 8645 438 8661 472
rect 8561 400 8661 438
rect 8719 472 8819 488
rect 8719 438 8735 472
rect 8803 438 8819 472
rect 8719 400 8819 438
rect 8877 472 8977 488
rect 8877 438 8893 472
rect 8961 438 8977 472
rect 8877 400 8977 438
rect 9035 472 9135 488
rect 9035 438 9051 472
rect 9119 438 9135 472
rect 9035 400 9135 438
rect 9193 472 9293 488
rect 9193 438 9209 472
rect 9277 438 9293 472
rect 9193 400 9293 438
rect 9351 472 9451 488
rect 9351 438 9367 472
rect 9435 438 9451 472
rect 9351 400 9451 438
rect 9509 472 9609 488
rect 9509 438 9525 472
rect 9593 438 9609 472
rect 9509 400 9609 438
rect 9667 472 9767 488
rect 9667 438 9683 472
rect 9751 438 9767 472
rect 9667 400 9767 438
rect 9825 472 9925 488
rect 9825 438 9841 472
rect 9909 438 9925 472
rect 9825 400 9925 438
rect 9983 472 10083 488
rect 9983 438 9999 472
rect 10067 438 10083 472
rect 9983 400 10083 438
rect 10141 472 10241 488
rect 10141 438 10157 472
rect 10225 438 10241 472
rect 10141 400 10241 438
rect 10299 472 10399 488
rect 10299 438 10315 472
rect 10383 438 10399 472
rect 10299 400 10399 438
rect 10457 472 10557 488
rect 10457 438 10473 472
rect 10541 438 10557 472
rect 10457 400 10557 438
rect 10615 472 10715 488
rect 10615 438 10631 472
rect 10699 438 10715 472
rect 10615 400 10715 438
rect 10773 472 10873 488
rect 10773 438 10789 472
rect 10857 438 10873 472
rect 10773 400 10873 438
rect 10931 472 11031 488
rect 10931 438 10947 472
rect 11015 438 11031 472
rect 10931 400 11031 438
rect 11089 472 11189 488
rect 11089 438 11105 472
rect 11173 438 11189 472
rect 11089 400 11189 438
rect 11247 472 11347 488
rect 11247 438 11263 472
rect 11331 438 11347 472
rect 11247 400 11347 438
rect 11405 472 11505 488
rect 11405 438 11421 472
rect 11489 438 11505 472
rect 11405 400 11505 438
rect 11563 472 11663 488
rect 11563 438 11579 472
rect 11647 438 11663 472
rect 11563 400 11663 438
rect 11721 472 11821 488
rect 11721 438 11737 472
rect 11805 438 11821 472
rect 11721 400 11821 438
rect 11879 472 11979 488
rect 11879 438 11895 472
rect 11963 438 11979 472
rect 11879 400 11979 438
rect 12037 472 12137 488
rect 12037 438 12053 472
rect 12121 438 12137 472
rect 12037 400 12137 438
rect 12195 472 12295 488
rect 12195 438 12211 472
rect 12279 438 12295 472
rect 12195 400 12295 438
rect 12353 472 12453 488
rect 12353 438 12369 472
rect 12437 438 12453 472
rect 12353 400 12453 438
rect 12511 472 12611 488
rect 12511 438 12527 472
rect 12595 438 12611 472
rect 12511 400 12611 438
rect 12669 472 12769 488
rect 12669 438 12685 472
rect 12753 438 12769 472
rect 12669 400 12769 438
rect 12827 472 12927 488
rect 12827 438 12843 472
rect 12911 438 12927 472
rect 12827 400 12927 438
rect -12927 -438 -12827 -400
rect -12927 -472 -12911 -438
rect -12843 -472 -12827 -438
rect -12927 -488 -12827 -472
rect -12769 -438 -12669 -400
rect -12769 -472 -12753 -438
rect -12685 -472 -12669 -438
rect -12769 -488 -12669 -472
rect -12611 -438 -12511 -400
rect -12611 -472 -12595 -438
rect -12527 -472 -12511 -438
rect -12611 -488 -12511 -472
rect -12453 -438 -12353 -400
rect -12453 -472 -12437 -438
rect -12369 -472 -12353 -438
rect -12453 -488 -12353 -472
rect -12295 -438 -12195 -400
rect -12295 -472 -12279 -438
rect -12211 -472 -12195 -438
rect -12295 -488 -12195 -472
rect -12137 -438 -12037 -400
rect -12137 -472 -12121 -438
rect -12053 -472 -12037 -438
rect -12137 -488 -12037 -472
rect -11979 -438 -11879 -400
rect -11979 -472 -11963 -438
rect -11895 -472 -11879 -438
rect -11979 -488 -11879 -472
rect -11821 -438 -11721 -400
rect -11821 -472 -11805 -438
rect -11737 -472 -11721 -438
rect -11821 -488 -11721 -472
rect -11663 -438 -11563 -400
rect -11663 -472 -11647 -438
rect -11579 -472 -11563 -438
rect -11663 -488 -11563 -472
rect -11505 -438 -11405 -400
rect -11505 -472 -11489 -438
rect -11421 -472 -11405 -438
rect -11505 -488 -11405 -472
rect -11347 -438 -11247 -400
rect -11347 -472 -11331 -438
rect -11263 -472 -11247 -438
rect -11347 -488 -11247 -472
rect -11189 -438 -11089 -400
rect -11189 -472 -11173 -438
rect -11105 -472 -11089 -438
rect -11189 -488 -11089 -472
rect -11031 -438 -10931 -400
rect -11031 -472 -11015 -438
rect -10947 -472 -10931 -438
rect -11031 -488 -10931 -472
rect -10873 -438 -10773 -400
rect -10873 -472 -10857 -438
rect -10789 -472 -10773 -438
rect -10873 -488 -10773 -472
rect -10715 -438 -10615 -400
rect -10715 -472 -10699 -438
rect -10631 -472 -10615 -438
rect -10715 -488 -10615 -472
rect -10557 -438 -10457 -400
rect -10557 -472 -10541 -438
rect -10473 -472 -10457 -438
rect -10557 -488 -10457 -472
rect -10399 -438 -10299 -400
rect -10399 -472 -10383 -438
rect -10315 -472 -10299 -438
rect -10399 -488 -10299 -472
rect -10241 -438 -10141 -400
rect -10241 -472 -10225 -438
rect -10157 -472 -10141 -438
rect -10241 -488 -10141 -472
rect -10083 -438 -9983 -400
rect -10083 -472 -10067 -438
rect -9999 -472 -9983 -438
rect -10083 -488 -9983 -472
rect -9925 -438 -9825 -400
rect -9925 -472 -9909 -438
rect -9841 -472 -9825 -438
rect -9925 -488 -9825 -472
rect -9767 -438 -9667 -400
rect -9767 -472 -9751 -438
rect -9683 -472 -9667 -438
rect -9767 -488 -9667 -472
rect -9609 -438 -9509 -400
rect -9609 -472 -9593 -438
rect -9525 -472 -9509 -438
rect -9609 -488 -9509 -472
rect -9451 -438 -9351 -400
rect -9451 -472 -9435 -438
rect -9367 -472 -9351 -438
rect -9451 -488 -9351 -472
rect -9293 -438 -9193 -400
rect -9293 -472 -9277 -438
rect -9209 -472 -9193 -438
rect -9293 -488 -9193 -472
rect -9135 -438 -9035 -400
rect -9135 -472 -9119 -438
rect -9051 -472 -9035 -438
rect -9135 -488 -9035 -472
rect -8977 -438 -8877 -400
rect -8977 -472 -8961 -438
rect -8893 -472 -8877 -438
rect -8977 -488 -8877 -472
rect -8819 -438 -8719 -400
rect -8819 -472 -8803 -438
rect -8735 -472 -8719 -438
rect -8819 -488 -8719 -472
rect -8661 -438 -8561 -400
rect -8661 -472 -8645 -438
rect -8577 -472 -8561 -438
rect -8661 -488 -8561 -472
rect -8503 -438 -8403 -400
rect -8503 -472 -8487 -438
rect -8419 -472 -8403 -438
rect -8503 -488 -8403 -472
rect -8345 -438 -8245 -400
rect -8345 -472 -8329 -438
rect -8261 -472 -8245 -438
rect -8345 -488 -8245 -472
rect -8187 -438 -8087 -400
rect -8187 -472 -8171 -438
rect -8103 -472 -8087 -438
rect -8187 -488 -8087 -472
rect -8029 -438 -7929 -400
rect -8029 -472 -8013 -438
rect -7945 -472 -7929 -438
rect -8029 -488 -7929 -472
rect -7871 -438 -7771 -400
rect -7871 -472 -7855 -438
rect -7787 -472 -7771 -438
rect -7871 -488 -7771 -472
rect -7713 -438 -7613 -400
rect -7713 -472 -7697 -438
rect -7629 -472 -7613 -438
rect -7713 -488 -7613 -472
rect -7555 -438 -7455 -400
rect -7555 -472 -7539 -438
rect -7471 -472 -7455 -438
rect -7555 -488 -7455 -472
rect -7397 -438 -7297 -400
rect -7397 -472 -7381 -438
rect -7313 -472 -7297 -438
rect -7397 -488 -7297 -472
rect -7239 -438 -7139 -400
rect -7239 -472 -7223 -438
rect -7155 -472 -7139 -438
rect -7239 -488 -7139 -472
rect -7081 -438 -6981 -400
rect -7081 -472 -7065 -438
rect -6997 -472 -6981 -438
rect -7081 -488 -6981 -472
rect -6923 -438 -6823 -400
rect -6923 -472 -6907 -438
rect -6839 -472 -6823 -438
rect -6923 -488 -6823 -472
rect -6765 -438 -6665 -400
rect -6765 -472 -6749 -438
rect -6681 -472 -6665 -438
rect -6765 -488 -6665 -472
rect -6607 -438 -6507 -400
rect -6607 -472 -6591 -438
rect -6523 -472 -6507 -438
rect -6607 -488 -6507 -472
rect -6449 -438 -6349 -400
rect -6449 -472 -6433 -438
rect -6365 -472 -6349 -438
rect -6449 -488 -6349 -472
rect -6291 -438 -6191 -400
rect -6291 -472 -6275 -438
rect -6207 -472 -6191 -438
rect -6291 -488 -6191 -472
rect -6133 -438 -6033 -400
rect -6133 -472 -6117 -438
rect -6049 -472 -6033 -438
rect -6133 -488 -6033 -472
rect -5975 -438 -5875 -400
rect -5975 -472 -5959 -438
rect -5891 -472 -5875 -438
rect -5975 -488 -5875 -472
rect -5817 -438 -5717 -400
rect -5817 -472 -5801 -438
rect -5733 -472 -5717 -438
rect -5817 -488 -5717 -472
rect -5659 -438 -5559 -400
rect -5659 -472 -5643 -438
rect -5575 -472 -5559 -438
rect -5659 -488 -5559 -472
rect -5501 -438 -5401 -400
rect -5501 -472 -5485 -438
rect -5417 -472 -5401 -438
rect -5501 -488 -5401 -472
rect -5343 -438 -5243 -400
rect -5343 -472 -5327 -438
rect -5259 -472 -5243 -438
rect -5343 -488 -5243 -472
rect -5185 -438 -5085 -400
rect -5185 -472 -5169 -438
rect -5101 -472 -5085 -438
rect -5185 -488 -5085 -472
rect -5027 -438 -4927 -400
rect -5027 -472 -5011 -438
rect -4943 -472 -4927 -438
rect -5027 -488 -4927 -472
rect -4869 -438 -4769 -400
rect -4869 -472 -4853 -438
rect -4785 -472 -4769 -438
rect -4869 -488 -4769 -472
rect -4711 -438 -4611 -400
rect -4711 -472 -4695 -438
rect -4627 -472 -4611 -438
rect -4711 -488 -4611 -472
rect -4553 -438 -4453 -400
rect -4553 -472 -4537 -438
rect -4469 -472 -4453 -438
rect -4553 -488 -4453 -472
rect -4395 -438 -4295 -400
rect -4395 -472 -4379 -438
rect -4311 -472 -4295 -438
rect -4395 -488 -4295 -472
rect -4237 -438 -4137 -400
rect -4237 -472 -4221 -438
rect -4153 -472 -4137 -438
rect -4237 -488 -4137 -472
rect -4079 -438 -3979 -400
rect -4079 -472 -4063 -438
rect -3995 -472 -3979 -438
rect -4079 -488 -3979 -472
rect -3921 -438 -3821 -400
rect -3921 -472 -3905 -438
rect -3837 -472 -3821 -438
rect -3921 -488 -3821 -472
rect -3763 -438 -3663 -400
rect -3763 -472 -3747 -438
rect -3679 -472 -3663 -438
rect -3763 -488 -3663 -472
rect -3605 -438 -3505 -400
rect -3605 -472 -3589 -438
rect -3521 -472 -3505 -438
rect -3605 -488 -3505 -472
rect -3447 -438 -3347 -400
rect -3447 -472 -3431 -438
rect -3363 -472 -3347 -438
rect -3447 -488 -3347 -472
rect -3289 -438 -3189 -400
rect -3289 -472 -3273 -438
rect -3205 -472 -3189 -438
rect -3289 -488 -3189 -472
rect -3131 -438 -3031 -400
rect -3131 -472 -3115 -438
rect -3047 -472 -3031 -438
rect -3131 -488 -3031 -472
rect -2973 -438 -2873 -400
rect -2973 -472 -2957 -438
rect -2889 -472 -2873 -438
rect -2973 -488 -2873 -472
rect -2815 -438 -2715 -400
rect -2815 -472 -2799 -438
rect -2731 -472 -2715 -438
rect -2815 -488 -2715 -472
rect -2657 -438 -2557 -400
rect -2657 -472 -2641 -438
rect -2573 -472 -2557 -438
rect -2657 -488 -2557 -472
rect -2499 -438 -2399 -400
rect -2499 -472 -2483 -438
rect -2415 -472 -2399 -438
rect -2499 -488 -2399 -472
rect -2341 -438 -2241 -400
rect -2341 -472 -2325 -438
rect -2257 -472 -2241 -438
rect -2341 -488 -2241 -472
rect -2183 -438 -2083 -400
rect -2183 -472 -2167 -438
rect -2099 -472 -2083 -438
rect -2183 -488 -2083 -472
rect -2025 -438 -1925 -400
rect -2025 -472 -2009 -438
rect -1941 -472 -1925 -438
rect -2025 -488 -1925 -472
rect -1867 -438 -1767 -400
rect -1867 -472 -1851 -438
rect -1783 -472 -1767 -438
rect -1867 -488 -1767 -472
rect -1709 -438 -1609 -400
rect -1709 -472 -1693 -438
rect -1625 -472 -1609 -438
rect -1709 -488 -1609 -472
rect -1551 -438 -1451 -400
rect -1551 -472 -1535 -438
rect -1467 -472 -1451 -438
rect -1551 -488 -1451 -472
rect -1393 -438 -1293 -400
rect -1393 -472 -1377 -438
rect -1309 -472 -1293 -438
rect -1393 -488 -1293 -472
rect -1235 -438 -1135 -400
rect -1235 -472 -1219 -438
rect -1151 -472 -1135 -438
rect -1235 -488 -1135 -472
rect -1077 -438 -977 -400
rect -1077 -472 -1061 -438
rect -993 -472 -977 -438
rect -1077 -488 -977 -472
rect -919 -438 -819 -400
rect -919 -472 -903 -438
rect -835 -472 -819 -438
rect -919 -488 -819 -472
rect -761 -438 -661 -400
rect -761 -472 -745 -438
rect -677 -472 -661 -438
rect -761 -488 -661 -472
rect -603 -438 -503 -400
rect -603 -472 -587 -438
rect -519 -472 -503 -438
rect -603 -488 -503 -472
rect -445 -438 -345 -400
rect -445 -472 -429 -438
rect -361 -472 -345 -438
rect -445 -488 -345 -472
rect -287 -438 -187 -400
rect -287 -472 -271 -438
rect -203 -472 -187 -438
rect -287 -488 -187 -472
rect -129 -438 -29 -400
rect -129 -472 -113 -438
rect -45 -472 -29 -438
rect -129 -488 -29 -472
rect 29 -438 129 -400
rect 29 -472 45 -438
rect 113 -472 129 -438
rect 29 -488 129 -472
rect 187 -438 287 -400
rect 187 -472 203 -438
rect 271 -472 287 -438
rect 187 -488 287 -472
rect 345 -438 445 -400
rect 345 -472 361 -438
rect 429 -472 445 -438
rect 345 -488 445 -472
rect 503 -438 603 -400
rect 503 -472 519 -438
rect 587 -472 603 -438
rect 503 -488 603 -472
rect 661 -438 761 -400
rect 661 -472 677 -438
rect 745 -472 761 -438
rect 661 -488 761 -472
rect 819 -438 919 -400
rect 819 -472 835 -438
rect 903 -472 919 -438
rect 819 -488 919 -472
rect 977 -438 1077 -400
rect 977 -472 993 -438
rect 1061 -472 1077 -438
rect 977 -488 1077 -472
rect 1135 -438 1235 -400
rect 1135 -472 1151 -438
rect 1219 -472 1235 -438
rect 1135 -488 1235 -472
rect 1293 -438 1393 -400
rect 1293 -472 1309 -438
rect 1377 -472 1393 -438
rect 1293 -488 1393 -472
rect 1451 -438 1551 -400
rect 1451 -472 1467 -438
rect 1535 -472 1551 -438
rect 1451 -488 1551 -472
rect 1609 -438 1709 -400
rect 1609 -472 1625 -438
rect 1693 -472 1709 -438
rect 1609 -488 1709 -472
rect 1767 -438 1867 -400
rect 1767 -472 1783 -438
rect 1851 -472 1867 -438
rect 1767 -488 1867 -472
rect 1925 -438 2025 -400
rect 1925 -472 1941 -438
rect 2009 -472 2025 -438
rect 1925 -488 2025 -472
rect 2083 -438 2183 -400
rect 2083 -472 2099 -438
rect 2167 -472 2183 -438
rect 2083 -488 2183 -472
rect 2241 -438 2341 -400
rect 2241 -472 2257 -438
rect 2325 -472 2341 -438
rect 2241 -488 2341 -472
rect 2399 -438 2499 -400
rect 2399 -472 2415 -438
rect 2483 -472 2499 -438
rect 2399 -488 2499 -472
rect 2557 -438 2657 -400
rect 2557 -472 2573 -438
rect 2641 -472 2657 -438
rect 2557 -488 2657 -472
rect 2715 -438 2815 -400
rect 2715 -472 2731 -438
rect 2799 -472 2815 -438
rect 2715 -488 2815 -472
rect 2873 -438 2973 -400
rect 2873 -472 2889 -438
rect 2957 -472 2973 -438
rect 2873 -488 2973 -472
rect 3031 -438 3131 -400
rect 3031 -472 3047 -438
rect 3115 -472 3131 -438
rect 3031 -488 3131 -472
rect 3189 -438 3289 -400
rect 3189 -472 3205 -438
rect 3273 -472 3289 -438
rect 3189 -488 3289 -472
rect 3347 -438 3447 -400
rect 3347 -472 3363 -438
rect 3431 -472 3447 -438
rect 3347 -488 3447 -472
rect 3505 -438 3605 -400
rect 3505 -472 3521 -438
rect 3589 -472 3605 -438
rect 3505 -488 3605 -472
rect 3663 -438 3763 -400
rect 3663 -472 3679 -438
rect 3747 -472 3763 -438
rect 3663 -488 3763 -472
rect 3821 -438 3921 -400
rect 3821 -472 3837 -438
rect 3905 -472 3921 -438
rect 3821 -488 3921 -472
rect 3979 -438 4079 -400
rect 3979 -472 3995 -438
rect 4063 -472 4079 -438
rect 3979 -488 4079 -472
rect 4137 -438 4237 -400
rect 4137 -472 4153 -438
rect 4221 -472 4237 -438
rect 4137 -488 4237 -472
rect 4295 -438 4395 -400
rect 4295 -472 4311 -438
rect 4379 -472 4395 -438
rect 4295 -488 4395 -472
rect 4453 -438 4553 -400
rect 4453 -472 4469 -438
rect 4537 -472 4553 -438
rect 4453 -488 4553 -472
rect 4611 -438 4711 -400
rect 4611 -472 4627 -438
rect 4695 -472 4711 -438
rect 4611 -488 4711 -472
rect 4769 -438 4869 -400
rect 4769 -472 4785 -438
rect 4853 -472 4869 -438
rect 4769 -488 4869 -472
rect 4927 -438 5027 -400
rect 4927 -472 4943 -438
rect 5011 -472 5027 -438
rect 4927 -488 5027 -472
rect 5085 -438 5185 -400
rect 5085 -472 5101 -438
rect 5169 -472 5185 -438
rect 5085 -488 5185 -472
rect 5243 -438 5343 -400
rect 5243 -472 5259 -438
rect 5327 -472 5343 -438
rect 5243 -488 5343 -472
rect 5401 -438 5501 -400
rect 5401 -472 5417 -438
rect 5485 -472 5501 -438
rect 5401 -488 5501 -472
rect 5559 -438 5659 -400
rect 5559 -472 5575 -438
rect 5643 -472 5659 -438
rect 5559 -488 5659 -472
rect 5717 -438 5817 -400
rect 5717 -472 5733 -438
rect 5801 -472 5817 -438
rect 5717 -488 5817 -472
rect 5875 -438 5975 -400
rect 5875 -472 5891 -438
rect 5959 -472 5975 -438
rect 5875 -488 5975 -472
rect 6033 -438 6133 -400
rect 6033 -472 6049 -438
rect 6117 -472 6133 -438
rect 6033 -488 6133 -472
rect 6191 -438 6291 -400
rect 6191 -472 6207 -438
rect 6275 -472 6291 -438
rect 6191 -488 6291 -472
rect 6349 -438 6449 -400
rect 6349 -472 6365 -438
rect 6433 -472 6449 -438
rect 6349 -488 6449 -472
rect 6507 -438 6607 -400
rect 6507 -472 6523 -438
rect 6591 -472 6607 -438
rect 6507 -488 6607 -472
rect 6665 -438 6765 -400
rect 6665 -472 6681 -438
rect 6749 -472 6765 -438
rect 6665 -488 6765 -472
rect 6823 -438 6923 -400
rect 6823 -472 6839 -438
rect 6907 -472 6923 -438
rect 6823 -488 6923 -472
rect 6981 -438 7081 -400
rect 6981 -472 6997 -438
rect 7065 -472 7081 -438
rect 6981 -488 7081 -472
rect 7139 -438 7239 -400
rect 7139 -472 7155 -438
rect 7223 -472 7239 -438
rect 7139 -488 7239 -472
rect 7297 -438 7397 -400
rect 7297 -472 7313 -438
rect 7381 -472 7397 -438
rect 7297 -488 7397 -472
rect 7455 -438 7555 -400
rect 7455 -472 7471 -438
rect 7539 -472 7555 -438
rect 7455 -488 7555 -472
rect 7613 -438 7713 -400
rect 7613 -472 7629 -438
rect 7697 -472 7713 -438
rect 7613 -488 7713 -472
rect 7771 -438 7871 -400
rect 7771 -472 7787 -438
rect 7855 -472 7871 -438
rect 7771 -488 7871 -472
rect 7929 -438 8029 -400
rect 7929 -472 7945 -438
rect 8013 -472 8029 -438
rect 7929 -488 8029 -472
rect 8087 -438 8187 -400
rect 8087 -472 8103 -438
rect 8171 -472 8187 -438
rect 8087 -488 8187 -472
rect 8245 -438 8345 -400
rect 8245 -472 8261 -438
rect 8329 -472 8345 -438
rect 8245 -488 8345 -472
rect 8403 -438 8503 -400
rect 8403 -472 8419 -438
rect 8487 -472 8503 -438
rect 8403 -488 8503 -472
rect 8561 -438 8661 -400
rect 8561 -472 8577 -438
rect 8645 -472 8661 -438
rect 8561 -488 8661 -472
rect 8719 -438 8819 -400
rect 8719 -472 8735 -438
rect 8803 -472 8819 -438
rect 8719 -488 8819 -472
rect 8877 -438 8977 -400
rect 8877 -472 8893 -438
rect 8961 -472 8977 -438
rect 8877 -488 8977 -472
rect 9035 -438 9135 -400
rect 9035 -472 9051 -438
rect 9119 -472 9135 -438
rect 9035 -488 9135 -472
rect 9193 -438 9293 -400
rect 9193 -472 9209 -438
rect 9277 -472 9293 -438
rect 9193 -488 9293 -472
rect 9351 -438 9451 -400
rect 9351 -472 9367 -438
rect 9435 -472 9451 -438
rect 9351 -488 9451 -472
rect 9509 -438 9609 -400
rect 9509 -472 9525 -438
rect 9593 -472 9609 -438
rect 9509 -488 9609 -472
rect 9667 -438 9767 -400
rect 9667 -472 9683 -438
rect 9751 -472 9767 -438
rect 9667 -488 9767 -472
rect 9825 -438 9925 -400
rect 9825 -472 9841 -438
rect 9909 -472 9925 -438
rect 9825 -488 9925 -472
rect 9983 -438 10083 -400
rect 9983 -472 9999 -438
rect 10067 -472 10083 -438
rect 9983 -488 10083 -472
rect 10141 -438 10241 -400
rect 10141 -472 10157 -438
rect 10225 -472 10241 -438
rect 10141 -488 10241 -472
rect 10299 -438 10399 -400
rect 10299 -472 10315 -438
rect 10383 -472 10399 -438
rect 10299 -488 10399 -472
rect 10457 -438 10557 -400
rect 10457 -472 10473 -438
rect 10541 -472 10557 -438
rect 10457 -488 10557 -472
rect 10615 -438 10715 -400
rect 10615 -472 10631 -438
rect 10699 -472 10715 -438
rect 10615 -488 10715 -472
rect 10773 -438 10873 -400
rect 10773 -472 10789 -438
rect 10857 -472 10873 -438
rect 10773 -488 10873 -472
rect 10931 -438 11031 -400
rect 10931 -472 10947 -438
rect 11015 -472 11031 -438
rect 10931 -488 11031 -472
rect 11089 -438 11189 -400
rect 11089 -472 11105 -438
rect 11173 -472 11189 -438
rect 11089 -488 11189 -472
rect 11247 -438 11347 -400
rect 11247 -472 11263 -438
rect 11331 -472 11347 -438
rect 11247 -488 11347 -472
rect 11405 -438 11505 -400
rect 11405 -472 11421 -438
rect 11489 -472 11505 -438
rect 11405 -488 11505 -472
rect 11563 -438 11663 -400
rect 11563 -472 11579 -438
rect 11647 -472 11663 -438
rect 11563 -488 11663 -472
rect 11721 -438 11821 -400
rect 11721 -472 11737 -438
rect 11805 -472 11821 -438
rect 11721 -488 11821 -472
rect 11879 -438 11979 -400
rect 11879 -472 11895 -438
rect 11963 -472 11979 -438
rect 11879 -488 11979 -472
rect 12037 -438 12137 -400
rect 12037 -472 12053 -438
rect 12121 -472 12137 -438
rect 12037 -488 12137 -472
rect 12195 -438 12295 -400
rect 12195 -472 12211 -438
rect 12279 -472 12295 -438
rect 12195 -488 12295 -472
rect 12353 -438 12453 -400
rect 12353 -472 12369 -438
rect 12437 -472 12453 -438
rect 12353 -488 12453 -472
rect 12511 -438 12611 -400
rect 12511 -472 12527 -438
rect 12595 -472 12611 -438
rect 12511 -488 12611 -472
rect 12669 -438 12769 -400
rect 12669 -472 12685 -438
rect 12753 -472 12769 -438
rect 12669 -488 12769 -472
rect 12827 -438 12927 -400
rect 12827 -472 12843 -438
rect 12911 -472 12927 -438
rect 12827 -488 12927 -472
<< polycont >>
rect -12911 438 -12843 472
rect -12753 438 -12685 472
rect -12595 438 -12527 472
rect -12437 438 -12369 472
rect -12279 438 -12211 472
rect -12121 438 -12053 472
rect -11963 438 -11895 472
rect -11805 438 -11737 472
rect -11647 438 -11579 472
rect -11489 438 -11421 472
rect -11331 438 -11263 472
rect -11173 438 -11105 472
rect -11015 438 -10947 472
rect -10857 438 -10789 472
rect -10699 438 -10631 472
rect -10541 438 -10473 472
rect -10383 438 -10315 472
rect -10225 438 -10157 472
rect -10067 438 -9999 472
rect -9909 438 -9841 472
rect -9751 438 -9683 472
rect -9593 438 -9525 472
rect -9435 438 -9367 472
rect -9277 438 -9209 472
rect -9119 438 -9051 472
rect -8961 438 -8893 472
rect -8803 438 -8735 472
rect -8645 438 -8577 472
rect -8487 438 -8419 472
rect -8329 438 -8261 472
rect -8171 438 -8103 472
rect -8013 438 -7945 472
rect -7855 438 -7787 472
rect -7697 438 -7629 472
rect -7539 438 -7471 472
rect -7381 438 -7313 472
rect -7223 438 -7155 472
rect -7065 438 -6997 472
rect -6907 438 -6839 472
rect -6749 438 -6681 472
rect -6591 438 -6523 472
rect -6433 438 -6365 472
rect -6275 438 -6207 472
rect -6117 438 -6049 472
rect -5959 438 -5891 472
rect -5801 438 -5733 472
rect -5643 438 -5575 472
rect -5485 438 -5417 472
rect -5327 438 -5259 472
rect -5169 438 -5101 472
rect -5011 438 -4943 472
rect -4853 438 -4785 472
rect -4695 438 -4627 472
rect -4537 438 -4469 472
rect -4379 438 -4311 472
rect -4221 438 -4153 472
rect -4063 438 -3995 472
rect -3905 438 -3837 472
rect -3747 438 -3679 472
rect -3589 438 -3521 472
rect -3431 438 -3363 472
rect -3273 438 -3205 472
rect -3115 438 -3047 472
rect -2957 438 -2889 472
rect -2799 438 -2731 472
rect -2641 438 -2573 472
rect -2483 438 -2415 472
rect -2325 438 -2257 472
rect -2167 438 -2099 472
rect -2009 438 -1941 472
rect -1851 438 -1783 472
rect -1693 438 -1625 472
rect -1535 438 -1467 472
rect -1377 438 -1309 472
rect -1219 438 -1151 472
rect -1061 438 -993 472
rect -903 438 -835 472
rect -745 438 -677 472
rect -587 438 -519 472
rect -429 438 -361 472
rect -271 438 -203 472
rect -113 438 -45 472
rect 45 438 113 472
rect 203 438 271 472
rect 361 438 429 472
rect 519 438 587 472
rect 677 438 745 472
rect 835 438 903 472
rect 993 438 1061 472
rect 1151 438 1219 472
rect 1309 438 1377 472
rect 1467 438 1535 472
rect 1625 438 1693 472
rect 1783 438 1851 472
rect 1941 438 2009 472
rect 2099 438 2167 472
rect 2257 438 2325 472
rect 2415 438 2483 472
rect 2573 438 2641 472
rect 2731 438 2799 472
rect 2889 438 2957 472
rect 3047 438 3115 472
rect 3205 438 3273 472
rect 3363 438 3431 472
rect 3521 438 3589 472
rect 3679 438 3747 472
rect 3837 438 3905 472
rect 3995 438 4063 472
rect 4153 438 4221 472
rect 4311 438 4379 472
rect 4469 438 4537 472
rect 4627 438 4695 472
rect 4785 438 4853 472
rect 4943 438 5011 472
rect 5101 438 5169 472
rect 5259 438 5327 472
rect 5417 438 5485 472
rect 5575 438 5643 472
rect 5733 438 5801 472
rect 5891 438 5959 472
rect 6049 438 6117 472
rect 6207 438 6275 472
rect 6365 438 6433 472
rect 6523 438 6591 472
rect 6681 438 6749 472
rect 6839 438 6907 472
rect 6997 438 7065 472
rect 7155 438 7223 472
rect 7313 438 7381 472
rect 7471 438 7539 472
rect 7629 438 7697 472
rect 7787 438 7855 472
rect 7945 438 8013 472
rect 8103 438 8171 472
rect 8261 438 8329 472
rect 8419 438 8487 472
rect 8577 438 8645 472
rect 8735 438 8803 472
rect 8893 438 8961 472
rect 9051 438 9119 472
rect 9209 438 9277 472
rect 9367 438 9435 472
rect 9525 438 9593 472
rect 9683 438 9751 472
rect 9841 438 9909 472
rect 9999 438 10067 472
rect 10157 438 10225 472
rect 10315 438 10383 472
rect 10473 438 10541 472
rect 10631 438 10699 472
rect 10789 438 10857 472
rect 10947 438 11015 472
rect 11105 438 11173 472
rect 11263 438 11331 472
rect 11421 438 11489 472
rect 11579 438 11647 472
rect 11737 438 11805 472
rect 11895 438 11963 472
rect 12053 438 12121 472
rect 12211 438 12279 472
rect 12369 438 12437 472
rect 12527 438 12595 472
rect 12685 438 12753 472
rect 12843 438 12911 472
rect -12911 -472 -12843 -438
rect -12753 -472 -12685 -438
rect -12595 -472 -12527 -438
rect -12437 -472 -12369 -438
rect -12279 -472 -12211 -438
rect -12121 -472 -12053 -438
rect -11963 -472 -11895 -438
rect -11805 -472 -11737 -438
rect -11647 -472 -11579 -438
rect -11489 -472 -11421 -438
rect -11331 -472 -11263 -438
rect -11173 -472 -11105 -438
rect -11015 -472 -10947 -438
rect -10857 -472 -10789 -438
rect -10699 -472 -10631 -438
rect -10541 -472 -10473 -438
rect -10383 -472 -10315 -438
rect -10225 -472 -10157 -438
rect -10067 -472 -9999 -438
rect -9909 -472 -9841 -438
rect -9751 -472 -9683 -438
rect -9593 -472 -9525 -438
rect -9435 -472 -9367 -438
rect -9277 -472 -9209 -438
rect -9119 -472 -9051 -438
rect -8961 -472 -8893 -438
rect -8803 -472 -8735 -438
rect -8645 -472 -8577 -438
rect -8487 -472 -8419 -438
rect -8329 -472 -8261 -438
rect -8171 -472 -8103 -438
rect -8013 -472 -7945 -438
rect -7855 -472 -7787 -438
rect -7697 -472 -7629 -438
rect -7539 -472 -7471 -438
rect -7381 -472 -7313 -438
rect -7223 -472 -7155 -438
rect -7065 -472 -6997 -438
rect -6907 -472 -6839 -438
rect -6749 -472 -6681 -438
rect -6591 -472 -6523 -438
rect -6433 -472 -6365 -438
rect -6275 -472 -6207 -438
rect -6117 -472 -6049 -438
rect -5959 -472 -5891 -438
rect -5801 -472 -5733 -438
rect -5643 -472 -5575 -438
rect -5485 -472 -5417 -438
rect -5327 -472 -5259 -438
rect -5169 -472 -5101 -438
rect -5011 -472 -4943 -438
rect -4853 -472 -4785 -438
rect -4695 -472 -4627 -438
rect -4537 -472 -4469 -438
rect -4379 -472 -4311 -438
rect -4221 -472 -4153 -438
rect -4063 -472 -3995 -438
rect -3905 -472 -3837 -438
rect -3747 -472 -3679 -438
rect -3589 -472 -3521 -438
rect -3431 -472 -3363 -438
rect -3273 -472 -3205 -438
rect -3115 -472 -3047 -438
rect -2957 -472 -2889 -438
rect -2799 -472 -2731 -438
rect -2641 -472 -2573 -438
rect -2483 -472 -2415 -438
rect -2325 -472 -2257 -438
rect -2167 -472 -2099 -438
rect -2009 -472 -1941 -438
rect -1851 -472 -1783 -438
rect -1693 -472 -1625 -438
rect -1535 -472 -1467 -438
rect -1377 -472 -1309 -438
rect -1219 -472 -1151 -438
rect -1061 -472 -993 -438
rect -903 -472 -835 -438
rect -745 -472 -677 -438
rect -587 -472 -519 -438
rect -429 -472 -361 -438
rect -271 -472 -203 -438
rect -113 -472 -45 -438
rect 45 -472 113 -438
rect 203 -472 271 -438
rect 361 -472 429 -438
rect 519 -472 587 -438
rect 677 -472 745 -438
rect 835 -472 903 -438
rect 993 -472 1061 -438
rect 1151 -472 1219 -438
rect 1309 -472 1377 -438
rect 1467 -472 1535 -438
rect 1625 -472 1693 -438
rect 1783 -472 1851 -438
rect 1941 -472 2009 -438
rect 2099 -472 2167 -438
rect 2257 -472 2325 -438
rect 2415 -472 2483 -438
rect 2573 -472 2641 -438
rect 2731 -472 2799 -438
rect 2889 -472 2957 -438
rect 3047 -472 3115 -438
rect 3205 -472 3273 -438
rect 3363 -472 3431 -438
rect 3521 -472 3589 -438
rect 3679 -472 3747 -438
rect 3837 -472 3905 -438
rect 3995 -472 4063 -438
rect 4153 -472 4221 -438
rect 4311 -472 4379 -438
rect 4469 -472 4537 -438
rect 4627 -472 4695 -438
rect 4785 -472 4853 -438
rect 4943 -472 5011 -438
rect 5101 -472 5169 -438
rect 5259 -472 5327 -438
rect 5417 -472 5485 -438
rect 5575 -472 5643 -438
rect 5733 -472 5801 -438
rect 5891 -472 5959 -438
rect 6049 -472 6117 -438
rect 6207 -472 6275 -438
rect 6365 -472 6433 -438
rect 6523 -472 6591 -438
rect 6681 -472 6749 -438
rect 6839 -472 6907 -438
rect 6997 -472 7065 -438
rect 7155 -472 7223 -438
rect 7313 -472 7381 -438
rect 7471 -472 7539 -438
rect 7629 -472 7697 -438
rect 7787 -472 7855 -438
rect 7945 -472 8013 -438
rect 8103 -472 8171 -438
rect 8261 -472 8329 -438
rect 8419 -472 8487 -438
rect 8577 -472 8645 -438
rect 8735 -472 8803 -438
rect 8893 -472 8961 -438
rect 9051 -472 9119 -438
rect 9209 -472 9277 -438
rect 9367 -472 9435 -438
rect 9525 -472 9593 -438
rect 9683 -472 9751 -438
rect 9841 -472 9909 -438
rect 9999 -472 10067 -438
rect 10157 -472 10225 -438
rect 10315 -472 10383 -438
rect 10473 -472 10541 -438
rect 10631 -472 10699 -438
rect 10789 -472 10857 -438
rect 10947 -472 11015 -438
rect 11105 -472 11173 -438
rect 11263 -472 11331 -438
rect 11421 -472 11489 -438
rect 11579 -472 11647 -438
rect 11737 -472 11805 -438
rect 11895 -472 11963 -438
rect 12053 -472 12121 -438
rect 12211 -472 12279 -438
rect 12369 -472 12437 -438
rect 12527 -472 12595 -438
rect 12685 -472 12753 -438
rect 12843 -472 12911 -438
<< locali >>
rect -13107 514 -13073 576
rect 13073 514 13107 576
rect -12927 438 -12911 472
rect -12843 438 -12753 472
rect -12685 438 -12595 472
rect -12527 438 -12437 472
rect -12369 438 -12279 472
rect -12211 438 -12121 472
rect -12053 438 -11963 472
rect -11895 438 -11805 472
rect -11737 438 -11647 472
rect -11579 438 -11489 472
rect -11421 438 -11331 472
rect -11263 438 -11173 472
rect -11105 438 -11015 472
rect -10947 438 -10857 472
rect -10789 438 -10699 472
rect -10631 438 -10541 472
rect -10473 438 -10383 472
rect -10315 438 -10225 472
rect -10157 438 -10067 472
rect -9999 438 -9909 472
rect -9841 438 -9751 472
rect -9683 438 -9593 472
rect -9525 438 -9435 472
rect -9367 438 -9277 472
rect -9209 438 -9119 472
rect -9051 438 -8961 472
rect -8893 438 -8803 472
rect -8735 438 -8645 472
rect -8577 438 -8487 472
rect -8419 438 -8329 472
rect -8261 438 -8171 472
rect -8103 438 -8013 472
rect -7945 438 -7855 472
rect -7787 438 -7697 472
rect -7629 438 -7539 472
rect -7471 438 -7381 472
rect -7313 438 -7223 472
rect -7155 438 -7065 472
rect -6997 438 -6907 472
rect -6839 438 -6749 472
rect -6681 438 -6591 472
rect -6523 438 -6433 472
rect -6365 438 -6275 472
rect -6207 438 -6117 472
rect -6049 438 -5959 472
rect -5891 438 -5801 472
rect -5733 438 -5643 472
rect -5575 438 -5485 472
rect -5417 438 -5327 472
rect -5259 438 -5169 472
rect -5101 438 -5011 472
rect -4943 438 -4853 472
rect -4785 438 -4695 472
rect -4627 438 -4537 472
rect -4469 438 -4379 472
rect -4311 438 -4221 472
rect -4153 438 -4063 472
rect -3995 438 -3905 472
rect -3837 438 -3747 472
rect -3679 438 -3589 472
rect -3521 438 -3431 472
rect -3363 438 -3273 472
rect -3205 438 -3115 472
rect -3047 438 -2957 472
rect -2889 438 -2799 472
rect -2731 438 -2641 472
rect -2573 438 -2483 472
rect -2415 438 -2325 472
rect -2257 438 -2167 472
rect -2099 438 -2009 472
rect -1941 438 -1851 472
rect -1783 438 -1693 472
rect -1625 438 -1535 472
rect -1467 438 -1377 472
rect -1309 438 -1219 472
rect -1151 438 -1061 472
rect -993 438 -903 472
rect -835 438 -745 472
rect -677 438 -587 472
rect -519 438 -429 472
rect -361 438 -271 472
rect -203 438 -113 472
rect -45 438 45 472
rect 113 438 203 472
rect 271 438 361 472
rect 429 438 519 472
rect 587 438 677 472
rect 745 438 835 472
rect 903 438 993 472
rect 1061 438 1151 472
rect 1219 438 1309 472
rect 1377 438 1467 472
rect 1535 438 1625 472
rect 1693 438 1783 472
rect 1851 438 1941 472
rect 2009 438 2099 472
rect 2167 438 2257 472
rect 2325 438 2415 472
rect 2483 438 2573 472
rect 2641 438 2731 472
rect 2799 438 2889 472
rect 2957 438 3047 472
rect 3115 438 3205 472
rect 3273 438 3363 472
rect 3431 438 3521 472
rect 3589 438 3679 472
rect 3747 438 3837 472
rect 3905 438 3995 472
rect 4063 438 4153 472
rect 4221 438 4311 472
rect 4379 438 4469 472
rect 4537 438 4627 472
rect 4695 438 4785 472
rect 4853 438 4943 472
rect 5011 438 5101 472
rect 5169 438 5259 472
rect 5327 438 5417 472
rect 5485 438 5575 472
rect 5643 438 5733 472
rect 5801 438 5891 472
rect 5959 438 6049 472
rect 6117 438 6207 472
rect 6275 438 6365 472
rect 6433 438 6523 472
rect 6591 438 6681 472
rect 6749 438 6839 472
rect 6907 438 6997 472
rect 7065 438 7155 472
rect 7223 438 7313 472
rect 7381 438 7471 472
rect 7539 438 7629 472
rect 7697 438 7787 472
rect 7855 438 7945 472
rect 8013 438 8103 472
rect 8171 438 8261 472
rect 8329 438 8419 472
rect 8487 438 8577 472
rect 8645 438 8735 472
rect 8803 438 8893 472
rect 8961 438 9051 472
rect 9119 438 9209 472
rect 9277 438 9367 472
rect 9435 438 9525 472
rect 9593 438 9683 472
rect 9751 438 9841 472
rect 9909 438 9999 472
rect 10067 438 10157 472
rect 10225 438 10315 472
rect 10383 438 10473 472
rect 10541 438 10631 472
rect 10699 438 10789 472
rect 10857 438 10947 472
rect 11015 438 11105 472
rect 11173 438 11263 472
rect 11331 438 11421 472
rect 11489 438 11579 472
rect 11647 438 11737 472
rect 11805 438 11895 472
rect 11963 438 12053 472
rect 12121 438 12211 472
rect 12279 438 12369 472
rect 12437 438 12527 472
rect 12595 438 12685 472
rect 12753 438 12843 472
rect 12911 438 12927 472
rect -12973 388 -12939 404
rect -12973 -404 -12939 -388
rect -12815 388 -12781 404
rect -12815 -404 -12781 -388
rect -12657 388 -12623 404
rect -12657 -404 -12623 -388
rect -12499 388 -12465 404
rect -12499 -404 -12465 -388
rect -12341 388 -12307 404
rect -12341 -404 -12307 -388
rect -12183 388 -12149 404
rect -12183 -404 -12149 -388
rect -12025 388 -11991 404
rect -12025 -404 -11991 -388
rect -11867 388 -11833 404
rect -11867 -404 -11833 -388
rect -11709 388 -11675 404
rect -11709 -404 -11675 -388
rect -11551 388 -11517 404
rect -11551 -404 -11517 -388
rect -11393 388 -11359 404
rect -11393 -404 -11359 -388
rect -11235 388 -11201 404
rect -11235 -404 -11201 -388
rect -11077 388 -11043 404
rect -11077 -404 -11043 -388
rect -10919 388 -10885 404
rect -10919 -404 -10885 -388
rect -10761 388 -10727 404
rect -10761 -404 -10727 -388
rect -10603 388 -10569 404
rect -10603 -404 -10569 -388
rect -10445 388 -10411 404
rect -10445 -404 -10411 -388
rect -10287 388 -10253 404
rect -10287 -404 -10253 -388
rect -10129 388 -10095 404
rect -10129 -404 -10095 -388
rect -9971 388 -9937 404
rect -9971 -404 -9937 -388
rect -9813 388 -9779 404
rect -9813 -404 -9779 -388
rect -9655 388 -9621 404
rect -9655 -404 -9621 -388
rect -9497 388 -9463 404
rect -9497 -404 -9463 -388
rect -9339 388 -9305 404
rect -9339 -404 -9305 -388
rect -9181 388 -9147 404
rect -9181 -404 -9147 -388
rect -9023 388 -8989 404
rect -9023 -404 -8989 -388
rect -8865 388 -8831 404
rect -8865 -404 -8831 -388
rect -8707 388 -8673 404
rect -8707 -404 -8673 -388
rect -8549 388 -8515 404
rect -8549 -404 -8515 -388
rect -8391 388 -8357 404
rect -8391 -404 -8357 -388
rect -8233 388 -8199 404
rect -8233 -404 -8199 -388
rect -8075 388 -8041 404
rect -8075 -404 -8041 -388
rect -7917 388 -7883 404
rect -7917 -404 -7883 -388
rect -7759 388 -7725 404
rect -7759 -404 -7725 -388
rect -7601 388 -7567 404
rect -7601 -404 -7567 -388
rect -7443 388 -7409 404
rect -7443 -404 -7409 -388
rect -7285 388 -7251 404
rect -7285 -404 -7251 -388
rect -7127 388 -7093 404
rect -7127 -404 -7093 -388
rect -6969 388 -6935 404
rect -6969 -404 -6935 -388
rect -6811 388 -6777 404
rect -6811 -404 -6777 -388
rect -6653 388 -6619 404
rect -6653 -404 -6619 -388
rect -6495 388 -6461 404
rect -6495 -404 -6461 -388
rect -6337 388 -6303 404
rect -6337 -404 -6303 -388
rect -6179 388 -6145 404
rect -6179 -404 -6145 -388
rect -6021 388 -5987 404
rect -6021 -404 -5987 -388
rect -5863 388 -5829 404
rect -5863 -404 -5829 -388
rect -5705 388 -5671 404
rect -5705 -404 -5671 -388
rect -5547 388 -5513 404
rect -5547 -404 -5513 -388
rect -5389 388 -5355 404
rect -5389 -404 -5355 -388
rect -5231 388 -5197 404
rect -5231 -404 -5197 -388
rect -5073 388 -5039 404
rect -5073 -404 -5039 -388
rect -4915 388 -4881 404
rect -4915 -404 -4881 -388
rect -4757 388 -4723 404
rect -4757 -404 -4723 -388
rect -4599 388 -4565 438
rect -4599 -438 -4565 -388
rect -4441 388 -4407 404
rect -4441 -404 -4407 -388
rect -4283 388 -4249 404
rect -4283 -404 -4249 -388
rect -4125 388 -4091 404
rect -4125 -404 -4091 -388
rect -3967 388 -3933 404
rect -3967 -404 -3933 -388
rect -3809 388 -3775 404
rect -3809 -404 -3775 -388
rect -3651 388 -3617 404
rect -3651 -404 -3617 -388
rect -3493 388 -3459 404
rect -3493 -404 -3459 -388
rect -3335 388 -3301 404
rect -3335 -404 -3301 -388
rect -3177 388 -3143 404
rect -3177 -404 -3143 -388
rect -3019 388 -2985 404
rect -3019 -404 -2985 -388
rect -2861 388 -2827 404
rect -2861 -404 -2827 -388
rect -2703 388 -2669 404
rect -2703 -404 -2669 -388
rect -2545 388 -2511 404
rect -2545 -404 -2511 -388
rect -2387 388 -2353 404
rect -2387 -404 -2353 -388
rect -2229 388 -2195 404
rect -2229 -404 -2195 -388
rect -2071 388 -2037 404
rect -2071 -404 -2037 -388
rect -1913 388 -1879 404
rect -1913 -404 -1879 -388
rect -1755 388 -1721 404
rect -1755 -404 -1721 -388
rect -1597 388 -1563 404
rect -1597 -404 -1563 -388
rect -1439 388 -1405 404
rect -1439 -404 -1405 -388
rect -1281 388 -1247 404
rect -1281 -404 -1247 -388
rect -1123 388 -1089 404
rect -1123 -404 -1089 -388
rect -965 388 -931 404
rect -965 -404 -931 -388
rect -807 388 -773 404
rect -807 -404 -773 -388
rect -649 388 -615 404
rect -649 -404 -615 -388
rect -491 388 -457 404
rect -491 -404 -457 -388
rect -333 388 -299 404
rect -333 -404 -299 -388
rect -175 388 -141 404
rect -175 -404 -141 -388
rect -17 388 17 404
rect -17 -404 17 -388
rect 141 388 175 404
rect 141 -404 175 -388
rect 299 388 333 404
rect 299 -404 333 -388
rect 457 388 491 404
rect 457 -404 491 -388
rect 615 388 649 404
rect 615 -404 649 -388
rect 773 388 807 404
rect 773 -404 807 -388
rect 931 388 965 404
rect 931 -404 965 -388
rect 1089 388 1123 404
rect 1089 -404 1123 -388
rect 1247 388 1281 404
rect 1247 -404 1281 -388
rect 1405 388 1439 404
rect 1405 -404 1439 -388
rect 1563 388 1597 404
rect 1563 -404 1597 -388
rect 1721 388 1755 404
rect 1721 -404 1755 -388
rect 1879 388 1913 404
rect 1879 -404 1913 -388
rect 2037 388 2071 404
rect 2037 -404 2071 -388
rect 2195 388 2229 404
rect 2195 -404 2229 -388
rect 2353 388 2387 404
rect 2353 -404 2387 -388
rect 2511 388 2545 404
rect 2511 -404 2545 -388
rect 2669 388 2703 404
rect 2669 -404 2703 -388
rect 2827 388 2861 404
rect 2827 -404 2861 -388
rect 2985 388 3019 404
rect 2985 -404 3019 -388
rect 3143 388 3177 404
rect 3143 -404 3177 -388
rect 3301 388 3335 404
rect 3301 -404 3335 -388
rect 3459 388 3493 404
rect 3459 -404 3493 -388
rect 3617 388 3651 404
rect 3617 -404 3651 -388
rect 3775 388 3809 404
rect 3775 -404 3809 -388
rect 3933 388 3967 404
rect 3933 -404 3967 -388
rect 4091 388 4125 404
rect 4091 -404 4125 -388
rect 4249 388 4283 404
rect 4249 -404 4283 -388
rect 4407 388 4441 404
rect 4407 -404 4441 -388
rect 4565 388 4599 438
rect 4565 -438 4599 -388
rect 4723 388 4757 404
rect 4723 -404 4757 -388
rect 4881 388 4915 404
rect 4881 -404 4915 -388
rect 5039 388 5073 404
rect 5039 -404 5073 -388
rect 5197 388 5231 404
rect 5197 -404 5231 -388
rect 5355 388 5389 404
rect 5355 -404 5389 -388
rect 5513 388 5547 404
rect 5513 -404 5547 -388
rect 5671 388 5705 404
rect 5671 -404 5705 -388
rect 5829 388 5863 404
rect 5829 -404 5863 -388
rect 5987 388 6021 404
rect 5987 -404 6021 -388
rect 6145 388 6179 404
rect 6145 -404 6179 -388
rect 6303 388 6337 404
rect 6303 -404 6337 -388
rect 6461 388 6495 404
rect 6461 -404 6495 -388
rect 6619 388 6653 404
rect 6619 -404 6653 -388
rect 6777 388 6811 404
rect 6777 -404 6811 -388
rect 6935 388 6969 404
rect 6935 -404 6969 -388
rect 7093 388 7127 404
rect 7093 -404 7127 -388
rect 7251 388 7285 404
rect 7251 -404 7285 -388
rect 7409 388 7443 404
rect 7409 -404 7443 -388
rect 7567 388 7601 404
rect 7567 -404 7601 -388
rect 7725 388 7759 404
rect 7725 -404 7759 -388
rect 7883 388 7917 404
rect 7883 -404 7917 -388
rect 8041 388 8075 404
rect 8041 -404 8075 -388
rect 8199 388 8233 404
rect 8199 -404 8233 -388
rect 8357 388 8391 404
rect 8357 -404 8391 -388
rect 8515 388 8549 404
rect 8515 -404 8549 -388
rect 8673 388 8707 404
rect 8673 -404 8707 -388
rect 8831 388 8865 404
rect 8831 -404 8865 -388
rect 8989 388 9023 404
rect 8989 -404 9023 -388
rect 9147 388 9181 404
rect 9147 -404 9181 -388
rect 9305 388 9339 404
rect 9305 -404 9339 -388
rect 9463 388 9497 404
rect 9463 -404 9497 -388
rect 9621 388 9655 404
rect 9621 -404 9655 -388
rect 9779 388 9813 404
rect 9779 -404 9813 -388
rect 9937 388 9971 404
rect 9937 -404 9971 -388
rect 10095 388 10129 404
rect 10095 -404 10129 -388
rect 10253 388 10287 404
rect 10253 -404 10287 -388
rect 10411 388 10445 404
rect 10411 -404 10445 -388
rect 10569 388 10603 404
rect 10569 -404 10603 -388
rect 10727 388 10761 404
rect 10727 -404 10761 -388
rect 10885 388 10919 404
rect 10885 -404 10919 -388
rect 11043 388 11077 404
rect 11043 -404 11077 -388
rect 11201 388 11235 404
rect 11201 -404 11235 -388
rect 11359 388 11393 404
rect 11359 -404 11393 -388
rect 11517 388 11551 404
rect 11517 -404 11551 -388
rect 11675 388 11709 404
rect 11675 -404 11709 -388
rect 11833 388 11867 404
rect 11833 -404 11867 -388
rect 11991 388 12025 404
rect 11991 -404 12025 -388
rect 12149 388 12183 404
rect 12149 -404 12183 -388
rect 12307 388 12341 404
rect 12307 -404 12341 -388
rect 12465 388 12499 404
rect 12465 -404 12499 -388
rect 12623 388 12657 404
rect 12623 -404 12657 -388
rect 12781 388 12815 404
rect 12781 -404 12815 -388
rect 12939 388 12973 404
rect 12939 -404 12973 -388
rect -12927 -472 -12911 -438
rect -12843 -472 -12753 -438
rect -12685 -472 -12595 -438
rect -12527 -472 -12437 -438
rect -12369 -472 -12279 -438
rect -12211 -472 -12121 -438
rect -12053 -472 -11963 -438
rect -11895 -472 -11805 -438
rect -11737 -472 -11647 -438
rect -11579 -472 -11489 -438
rect -11421 -472 -11331 -438
rect -11263 -472 -11173 -438
rect -11105 -472 -11015 -438
rect -10947 -472 -10857 -438
rect -10789 -472 -10699 -438
rect -10631 -472 -10541 -438
rect -10473 -472 -10383 -438
rect -10315 -472 -10225 -438
rect -10157 -472 -10067 -438
rect -9999 -472 -9909 -438
rect -9841 -472 -9751 -438
rect -9683 -472 -9593 -438
rect -9525 -472 -9435 -438
rect -9367 -472 -9277 -438
rect -9209 -472 -9119 -438
rect -9051 -472 -8961 -438
rect -8893 -472 -8803 -438
rect -8735 -472 -8645 -438
rect -8577 -472 -8487 -438
rect -8419 -472 -8329 -438
rect -8261 -472 -8171 -438
rect -8103 -472 -8013 -438
rect -7945 -472 -7855 -438
rect -7787 -472 -7697 -438
rect -7629 -472 -7539 -438
rect -7471 -472 -7381 -438
rect -7313 -472 -7223 -438
rect -7155 -472 -7065 -438
rect -6997 -472 -6907 -438
rect -6839 -472 -6749 -438
rect -6681 -472 -6591 -438
rect -6523 -472 -6433 -438
rect -6365 -472 -6275 -438
rect -6207 -472 -6117 -438
rect -6049 -472 -5959 -438
rect -5891 -472 -5801 -438
rect -5733 -472 -5643 -438
rect -5575 -472 -5485 -438
rect -5417 -472 -5327 -438
rect -5259 -472 -5169 -438
rect -5101 -472 -5011 -438
rect -4943 -472 -4853 -438
rect -4785 -472 -4695 -438
rect -4627 -472 -4537 -438
rect -4469 -472 -4379 -438
rect -4311 -472 -4221 -438
rect -4153 -472 -4063 -438
rect -3995 -472 -3905 -438
rect -3837 -472 -3747 -438
rect -3679 -472 -3589 -438
rect -3521 -472 -3431 -438
rect -3363 -472 -3273 -438
rect -3205 -472 -3115 -438
rect -3047 -472 -2957 -438
rect -2889 -472 -2799 -438
rect -2731 -472 -2641 -438
rect -2573 -472 -2483 -438
rect -2415 -472 -2325 -438
rect -2257 -472 -2167 -438
rect -2099 -472 -2009 -438
rect -1941 -472 -1851 -438
rect -1783 -472 -1693 -438
rect -1625 -472 -1535 -438
rect -1467 -472 -1377 -438
rect -1309 -472 -1219 -438
rect -1151 -472 -1061 -438
rect -993 -472 -903 -438
rect -835 -472 -745 -438
rect -677 -472 -587 -438
rect -519 -472 -429 -438
rect -361 -472 -271 -438
rect -203 -472 -113 -438
rect -45 -472 45 -438
rect 113 -472 203 -438
rect 271 -472 361 -438
rect 429 -472 519 -438
rect 587 -472 677 -438
rect 745 -472 835 -438
rect 903 -472 993 -438
rect 1061 -472 1151 -438
rect 1219 -472 1309 -438
rect 1377 -472 1467 -438
rect 1535 -472 1625 -438
rect 1693 -472 1783 -438
rect 1851 -472 1941 -438
rect 2009 -472 2099 -438
rect 2167 -472 2257 -438
rect 2325 -472 2415 -438
rect 2483 -472 2573 -438
rect 2641 -472 2731 -438
rect 2799 -472 2889 -438
rect 2957 -472 3047 -438
rect 3115 -472 3205 -438
rect 3273 -472 3363 -438
rect 3431 -472 3521 -438
rect 3589 -472 3679 -438
rect 3747 -472 3837 -438
rect 3905 -472 3995 -438
rect 4063 -472 4153 -438
rect 4221 -472 4311 -438
rect 4379 -472 4469 -438
rect 4537 -472 4627 -438
rect 4695 -472 4785 -438
rect 4853 -472 4943 -438
rect 5011 -472 5101 -438
rect 5169 -472 5259 -438
rect 5327 -472 5417 -438
rect 5485 -472 5575 -438
rect 5643 -472 5733 -438
rect 5801 -472 5891 -438
rect 5959 -472 6049 -438
rect 6117 -472 6207 -438
rect 6275 -472 6365 -438
rect 6433 -472 6523 -438
rect 6591 -472 6681 -438
rect 6749 -472 6839 -438
rect 6907 -472 6997 -438
rect 7065 -472 7155 -438
rect 7223 -472 7313 -438
rect 7381 -472 7471 -438
rect 7539 -472 7629 -438
rect 7697 -472 7787 -438
rect 7855 -472 7945 -438
rect 8013 -472 8103 -438
rect 8171 -472 8261 -438
rect 8329 -472 8419 -438
rect 8487 -472 8577 -438
rect 8645 -472 8735 -438
rect 8803 -472 8893 -438
rect 8961 -472 9051 -438
rect 9119 -472 9209 -438
rect 9277 -472 9367 -438
rect 9435 -472 9525 -438
rect 9593 -472 9683 -438
rect 9751 -472 9841 -438
rect 9909 -472 9999 -438
rect 10067 -472 10157 -438
rect 10225 -472 10315 -438
rect 10383 -472 10473 -438
rect 10541 -472 10631 -438
rect 10699 -472 10789 -438
rect 10857 -472 10947 -438
rect 11015 -472 11105 -438
rect 11173 -472 11263 -438
rect 11331 -472 11421 -438
rect 11489 -472 11579 -438
rect 11647 -472 11737 -438
rect 11805 -472 11895 -438
rect 11963 -472 12053 -438
rect 12121 -472 12211 -438
rect 12279 -472 12369 -438
rect 12437 -472 12527 -438
rect 12595 -472 12685 -438
rect 12753 -472 12843 -438
rect 12911 -472 12927 -438
rect -13107 -576 -13073 -514
rect 13073 -576 13107 -514
<< viali >>
rect -13107 576 -13011 610
rect -13011 576 13011 610
rect 13011 576 13107 610
rect -12911 438 -12843 472
rect -12753 438 -12685 472
rect -12595 438 -12527 472
rect -12437 438 -12369 472
rect -12279 438 -12211 472
rect -12121 438 -12053 472
rect -11963 438 -11895 472
rect -11805 438 -11737 472
rect -11647 438 -11579 472
rect -11489 438 -11421 472
rect -11331 438 -11263 472
rect -11173 438 -11105 472
rect -11015 438 -10947 472
rect -10857 438 -10789 472
rect -10699 438 -10631 472
rect -10541 438 -10473 472
rect -10383 438 -10315 472
rect -10225 438 -10157 472
rect -10067 438 -9999 472
rect -9909 438 -9841 472
rect -9751 438 -9683 472
rect -9593 438 -9525 472
rect -9435 438 -9367 472
rect -9277 438 -9209 472
rect -9119 438 -9051 472
rect -8961 438 -8893 472
rect -8803 438 -8735 472
rect -8645 438 -8577 472
rect -8487 438 -8419 472
rect -8329 438 -8261 472
rect -8171 438 -8103 472
rect -8013 438 -7945 472
rect -7855 438 -7787 472
rect -7697 438 -7629 472
rect -7539 438 -7471 472
rect -7381 438 -7313 472
rect -7223 438 -7155 472
rect -7065 438 -6997 472
rect -6907 438 -6839 472
rect -6749 438 -6681 472
rect -6591 438 -6523 472
rect -6433 438 -6365 472
rect -6275 438 -6207 472
rect -6117 438 -6049 472
rect -5959 438 -5891 472
rect -5801 438 -5733 472
rect -5643 438 -5575 472
rect -5485 438 -5417 472
rect -5327 438 -5259 472
rect -5169 438 -5101 472
rect -5011 438 -4943 472
rect -4853 438 -4785 472
rect -4695 438 -4627 472
rect -4537 438 -4469 472
rect -4379 438 -4311 472
rect -4221 438 -4153 472
rect -4063 438 -3995 472
rect -3905 438 -3837 472
rect -3747 438 -3679 472
rect -3589 438 -3521 472
rect -3431 438 -3363 472
rect -3273 438 -3205 472
rect -3115 438 -3047 472
rect -2957 438 -2889 472
rect -2799 438 -2731 472
rect -2641 438 -2573 472
rect -2483 438 -2415 472
rect -2325 438 -2257 472
rect -2167 438 -2099 472
rect -2009 438 -1941 472
rect -1851 438 -1783 472
rect -1693 438 -1625 472
rect -1535 438 -1467 472
rect -1377 438 -1309 472
rect -1219 438 -1151 472
rect -1061 438 -993 472
rect -903 438 -835 472
rect -745 438 -677 472
rect -587 438 -519 472
rect -429 438 -361 472
rect -271 438 -203 472
rect -113 438 -45 472
rect 45 438 113 472
rect 203 438 271 472
rect 361 438 429 472
rect 519 438 587 472
rect 677 438 745 472
rect 835 438 903 472
rect 993 438 1061 472
rect 1151 438 1219 472
rect 1309 438 1377 472
rect 1467 438 1535 472
rect 1625 438 1693 472
rect 1783 438 1851 472
rect 1941 438 2009 472
rect 2099 438 2167 472
rect 2257 438 2325 472
rect 2415 438 2483 472
rect 2573 438 2641 472
rect 2731 438 2799 472
rect 2889 438 2957 472
rect 3047 438 3115 472
rect 3205 438 3273 472
rect 3363 438 3431 472
rect 3521 438 3589 472
rect 3679 438 3747 472
rect 3837 438 3905 472
rect 3995 438 4063 472
rect 4153 438 4221 472
rect 4311 438 4379 472
rect 4469 438 4537 472
rect 4627 438 4695 472
rect 4785 438 4853 472
rect 4943 438 5011 472
rect 5101 438 5169 472
rect 5259 438 5327 472
rect 5417 438 5485 472
rect 5575 438 5643 472
rect 5733 438 5801 472
rect 5891 438 5959 472
rect 6049 438 6117 472
rect 6207 438 6275 472
rect 6365 438 6433 472
rect 6523 438 6591 472
rect 6681 438 6749 472
rect 6839 438 6907 472
rect 6997 438 7065 472
rect 7155 438 7223 472
rect 7313 438 7381 472
rect 7471 438 7539 472
rect 7629 438 7697 472
rect 7787 438 7855 472
rect 7945 438 8013 472
rect 8103 438 8171 472
rect 8261 438 8329 472
rect 8419 438 8487 472
rect 8577 438 8645 472
rect 8735 438 8803 472
rect 8893 438 8961 472
rect 9051 438 9119 472
rect 9209 438 9277 472
rect 9367 438 9435 472
rect 9525 438 9593 472
rect 9683 438 9751 472
rect 9841 438 9909 472
rect 9999 438 10067 472
rect 10157 438 10225 472
rect 10315 438 10383 472
rect 10473 438 10541 472
rect 10631 438 10699 472
rect 10789 438 10857 472
rect 10947 438 11015 472
rect 11105 438 11173 472
rect 11263 438 11331 472
rect 11421 438 11489 472
rect 11579 438 11647 472
rect 11737 438 11805 472
rect 11895 438 11963 472
rect 12053 438 12121 472
rect 12211 438 12279 472
rect 12369 438 12437 472
rect 12527 438 12595 472
rect 12685 438 12753 472
rect 12843 438 12911 472
rect -12973 -388 -12939 388
rect -12815 -388 -12781 388
rect -12657 -388 -12623 388
rect -12499 -388 -12465 388
rect -12341 -388 -12307 388
rect -12183 -388 -12149 388
rect -12025 -388 -11991 388
rect -11867 -388 -11833 388
rect -11709 -388 -11675 388
rect -11551 -388 -11517 388
rect -11393 -388 -11359 388
rect -11235 -388 -11201 388
rect -11077 -388 -11043 388
rect -10919 -388 -10885 388
rect -10761 -388 -10727 388
rect -10603 -388 -10569 388
rect -10445 -388 -10411 388
rect -10287 -388 -10253 388
rect -10129 -388 -10095 388
rect -9971 -388 -9937 388
rect -9813 -388 -9779 388
rect -9655 -388 -9621 388
rect -9497 -388 -9463 388
rect -9339 -388 -9305 388
rect -9181 -388 -9147 388
rect -9023 -388 -8989 388
rect -8865 -388 -8831 388
rect -8707 -388 -8673 388
rect -8549 -388 -8515 388
rect -8391 -388 -8357 388
rect -8233 -388 -8199 388
rect -8075 -388 -8041 388
rect -7917 -388 -7883 388
rect -7759 -388 -7725 388
rect -7601 -388 -7567 388
rect -7443 -388 -7409 388
rect -7285 -388 -7251 388
rect -7127 -388 -7093 388
rect -6969 -388 -6935 388
rect -6811 -388 -6777 388
rect -6653 -388 -6619 388
rect -6495 -388 -6461 388
rect -6337 -388 -6303 388
rect -6179 -388 -6145 388
rect -6021 -388 -5987 388
rect -5863 -388 -5829 388
rect -5705 -388 -5671 388
rect -5547 -388 -5513 388
rect -5389 -388 -5355 388
rect -5231 -388 -5197 388
rect -5073 -388 -5039 388
rect -4915 -388 -4881 388
rect -4757 -388 -4723 388
rect -4599 -388 -4565 388
rect -4441 -388 -4407 388
rect -4283 -388 -4249 388
rect -4125 -388 -4091 388
rect -3967 -388 -3933 388
rect -3809 -388 -3775 388
rect -3651 -388 -3617 388
rect -3493 -388 -3459 388
rect -3335 -388 -3301 388
rect -3177 -388 -3143 388
rect -3019 -388 -2985 388
rect -2861 -388 -2827 388
rect -2703 -388 -2669 388
rect -2545 -388 -2511 388
rect -2387 -388 -2353 388
rect -2229 -388 -2195 388
rect -2071 -388 -2037 388
rect -1913 -388 -1879 388
rect -1755 -388 -1721 388
rect -1597 -388 -1563 388
rect -1439 -388 -1405 388
rect -1281 -388 -1247 388
rect -1123 -388 -1089 388
rect -965 -388 -931 388
rect -807 -388 -773 388
rect -649 -388 -615 388
rect -491 -388 -457 388
rect -333 -388 -299 388
rect -175 -388 -141 388
rect -17 -388 17 388
rect 141 -388 175 388
rect 299 -388 333 388
rect 457 -388 491 388
rect 615 -388 649 388
rect 773 -388 807 388
rect 931 -388 965 388
rect 1089 -388 1123 388
rect 1247 -388 1281 388
rect 1405 -388 1439 388
rect 1563 -388 1597 388
rect 1721 -388 1755 388
rect 1879 -388 1913 388
rect 2037 -388 2071 388
rect 2195 -388 2229 388
rect 2353 -388 2387 388
rect 2511 -388 2545 388
rect 2669 -388 2703 388
rect 2827 -388 2861 388
rect 2985 -388 3019 388
rect 3143 -388 3177 388
rect 3301 -388 3335 388
rect 3459 -388 3493 388
rect 3617 -388 3651 388
rect 3775 -388 3809 388
rect 3933 -388 3967 388
rect 4091 -388 4125 388
rect 4249 -388 4283 388
rect 4407 -388 4441 388
rect 4565 -388 4599 388
rect 4723 -388 4757 388
rect 4881 -388 4915 388
rect 5039 -388 5073 388
rect 5197 -388 5231 388
rect 5355 -388 5389 388
rect 5513 -388 5547 388
rect 5671 -388 5705 388
rect 5829 -388 5863 388
rect 5987 -388 6021 388
rect 6145 -388 6179 388
rect 6303 -388 6337 388
rect 6461 -388 6495 388
rect 6619 -388 6653 388
rect 6777 -388 6811 388
rect 6935 -388 6969 388
rect 7093 -388 7127 388
rect 7251 -388 7285 388
rect 7409 -388 7443 388
rect 7567 -388 7601 388
rect 7725 -388 7759 388
rect 7883 -388 7917 388
rect 8041 -388 8075 388
rect 8199 -388 8233 388
rect 8357 -388 8391 388
rect 8515 -388 8549 388
rect 8673 -388 8707 388
rect 8831 -388 8865 388
rect 8989 -388 9023 388
rect 9147 -388 9181 388
rect 9305 -388 9339 388
rect 9463 -388 9497 388
rect 9621 -388 9655 388
rect 9779 -388 9813 388
rect 9937 -388 9971 388
rect 10095 -388 10129 388
rect 10253 -388 10287 388
rect 10411 -388 10445 388
rect 10569 -388 10603 388
rect 10727 -388 10761 388
rect 10885 -388 10919 388
rect 11043 -388 11077 388
rect 11201 -388 11235 388
rect 11359 -388 11393 388
rect 11517 -388 11551 388
rect 11675 -388 11709 388
rect 11833 -388 11867 388
rect 11991 -388 12025 388
rect 12149 -388 12183 388
rect 12307 -388 12341 388
rect 12465 -388 12499 388
rect 12623 -388 12657 388
rect 12781 -388 12815 388
rect 12939 -388 12973 388
rect -12911 -472 -12843 -438
rect -12753 -472 -12685 -438
rect -12595 -472 -12527 -438
rect -12437 -472 -12369 -438
rect -12279 -472 -12211 -438
rect -12121 -472 -12053 -438
rect -11963 -472 -11895 -438
rect -11805 -472 -11737 -438
rect -11647 -472 -11579 -438
rect -11489 -472 -11421 -438
rect -11331 -472 -11263 -438
rect -11173 -472 -11105 -438
rect -11015 -472 -10947 -438
rect -10857 -472 -10789 -438
rect -10699 -472 -10631 -438
rect -10541 -472 -10473 -438
rect -10383 -472 -10315 -438
rect -10225 -472 -10157 -438
rect -10067 -472 -9999 -438
rect -9909 -472 -9841 -438
rect -9751 -472 -9683 -438
rect -9593 -472 -9525 -438
rect -9435 -472 -9367 -438
rect -9277 -472 -9209 -438
rect -9119 -472 -9051 -438
rect -8961 -472 -8893 -438
rect -8803 -472 -8735 -438
rect -8645 -472 -8577 -438
rect -8487 -472 -8419 -438
rect -8329 -472 -8261 -438
rect -8171 -472 -8103 -438
rect -8013 -472 -7945 -438
rect -7855 -472 -7787 -438
rect -7697 -472 -7629 -438
rect -7539 -472 -7471 -438
rect -7381 -472 -7313 -438
rect -7223 -472 -7155 -438
rect -7065 -472 -6997 -438
rect -6907 -472 -6839 -438
rect -6749 -472 -6681 -438
rect -6591 -472 -6523 -438
rect -6433 -472 -6365 -438
rect -6275 -472 -6207 -438
rect -6117 -472 -6049 -438
rect -5959 -472 -5891 -438
rect -5801 -472 -5733 -438
rect -5643 -472 -5575 -438
rect -5485 -472 -5417 -438
rect -5327 -472 -5259 -438
rect -5169 -472 -5101 -438
rect -5011 -472 -4943 -438
rect -4853 -472 -4785 -438
rect -4695 -472 -4627 -438
rect -4537 -472 -4469 -438
rect -4379 -472 -4311 -438
rect -4221 -472 -4153 -438
rect -4063 -472 -3995 -438
rect -3905 -472 -3837 -438
rect -3747 -472 -3679 -438
rect -3589 -472 -3521 -438
rect -3431 -472 -3363 -438
rect -3273 -472 -3205 -438
rect -3115 -472 -3047 -438
rect -2957 -472 -2889 -438
rect -2799 -472 -2731 -438
rect -2641 -472 -2573 -438
rect -2483 -472 -2415 -438
rect -2325 -472 -2257 -438
rect -2167 -472 -2099 -438
rect -2009 -472 -1941 -438
rect -1851 -472 -1783 -438
rect -1693 -472 -1625 -438
rect -1535 -472 -1467 -438
rect -1377 -472 -1309 -438
rect -1219 -472 -1151 -438
rect -1061 -472 -993 -438
rect -903 -472 -835 -438
rect -745 -472 -677 -438
rect -587 -472 -519 -438
rect -429 -472 -361 -438
rect -271 -472 -203 -438
rect -113 -472 -45 -438
rect 45 -472 113 -438
rect 203 -472 271 -438
rect 361 -472 429 -438
rect 519 -472 587 -438
rect 677 -472 745 -438
rect 835 -472 903 -438
rect 993 -472 1061 -438
rect 1151 -472 1219 -438
rect 1309 -472 1377 -438
rect 1467 -472 1535 -438
rect 1625 -472 1693 -438
rect 1783 -472 1851 -438
rect 1941 -472 2009 -438
rect 2099 -472 2167 -438
rect 2257 -472 2325 -438
rect 2415 -472 2483 -438
rect 2573 -472 2641 -438
rect 2731 -472 2799 -438
rect 2889 -472 2957 -438
rect 3047 -472 3115 -438
rect 3205 -472 3273 -438
rect 3363 -472 3431 -438
rect 3521 -472 3589 -438
rect 3679 -472 3747 -438
rect 3837 -472 3905 -438
rect 3995 -472 4063 -438
rect 4153 -472 4221 -438
rect 4311 -472 4379 -438
rect 4469 -472 4537 -438
rect 4627 -472 4695 -438
rect 4785 -472 4853 -438
rect 4943 -472 5011 -438
rect 5101 -472 5169 -438
rect 5259 -472 5327 -438
rect 5417 -472 5485 -438
rect 5575 -472 5643 -438
rect 5733 -472 5801 -438
rect 5891 -472 5959 -438
rect 6049 -472 6117 -438
rect 6207 -472 6275 -438
rect 6365 -472 6433 -438
rect 6523 -472 6591 -438
rect 6681 -472 6749 -438
rect 6839 -472 6907 -438
rect 6997 -472 7065 -438
rect 7155 -472 7223 -438
rect 7313 -472 7381 -438
rect 7471 -472 7539 -438
rect 7629 -472 7697 -438
rect 7787 -472 7855 -438
rect 7945 -472 8013 -438
rect 8103 -472 8171 -438
rect 8261 -472 8329 -438
rect 8419 -472 8487 -438
rect 8577 -472 8645 -438
rect 8735 -472 8803 -438
rect 8893 -472 8961 -438
rect 9051 -472 9119 -438
rect 9209 -472 9277 -438
rect 9367 -472 9435 -438
rect 9525 -472 9593 -438
rect 9683 -472 9751 -438
rect 9841 -472 9909 -438
rect 9999 -472 10067 -438
rect 10157 -472 10225 -438
rect 10315 -472 10383 -438
rect 10473 -472 10541 -438
rect 10631 -472 10699 -438
rect 10789 -472 10857 -438
rect 10947 -472 11015 -438
rect 11105 -472 11173 -438
rect 11263 -472 11331 -438
rect 11421 -472 11489 -438
rect 11579 -472 11647 -438
rect 11737 -472 11805 -438
rect 11895 -472 11963 -438
rect 12053 -472 12121 -438
rect 12211 -472 12279 -438
rect 12369 -472 12437 -438
rect 12527 -472 12595 -438
rect 12685 -472 12753 -438
rect 12843 -472 12911 -438
rect -13107 -610 -13011 -576
rect -13011 -610 13011 -576
rect 13011 -610 13107 -576
<< metal1 >>
rect -12990 616 -12984 619
rect -13119 610 -12984 616
rect -12928 616 -12922 619
rect -12674 616 -12668 619
rect -12928 610 -12668 616
rect -12612 616 -12606 619
rect -12358 616 -12352 619
rect -12612 610 -12352 616
rect -12296 616 -12290 619
rect -12042 616 -12036 619
rect -12296 610 -12036 616
rect -11980 616 -11974 619
rect -11726 616 -11720 619
rect -11980 610 -11720 616
rect -11664 616 -11658 619
rect -11410 616 -11404 619
rect -11664 610 -11404 616
rect -11348 616 -11342 619
rect -11094 616 -11088 619
rect -11348 610 -11088 616
rect -11032 616 -11026 619
rect -10778 616 -10772 619
rect -11032 610 -10772 616
rect -10716 616 -10710 619
rect -10462 616 -10456 619
rect -10716 610 -10456 616
rect -10400 616 -10394 619
rect -10146 616 -10140 619
rect -10400 610 -10140 616
rect -10084 616 -10078 619
rect -9830 616 -9824 619
rect -10084 610 -9824 616
rect -9768 616 -9762 619
rect -9514 616 -9508 619
rect -9768 610 -9508 616
rect -9452 616 -9446 619
rect -9198 616 -9192 619
rect -9452 610 -9192 616
rect -9136 616 -9130 619
rect -8882 616 -8876 619
rect -9136 610 -8876 616
rect -8820 616 -8814 619
rect -8566 616 -8560 619
rect -8820 610 -8560 616
rect -8504 616 -8498 619
rect -8250 616 -8244 619
rect -8504 610 -8244 616
rect -8188 616 -8182 619
rect -7934 616 -7928 619
rect -8188 610 -7928 616
rect -7872 616 -7866 619
rect -7618 616 -7612 619
rect -7872 610 -7612 616
rect -7556 616 -7550 619
rect -7302 616 -7296 619
rect -7556 610 -7296 616
rect -7240 616 -7234 619
rect -6986 616 -6980 619
rect -7240 610 -6980 616
rect -6924 616 -6918 619
rect -6670 616 -6664 619
rect -6924 610 -6664 616
rect -6608 616 -6602 619
rect -6354 616 -6348 619
rect -6608 610 -6348 616
rect -6292 616 -6286 619
rect -6038 616 -6032 619
rect -6292 610 -6032 616
rect -5976 616 -5970 619
rect -5722 616 -5716 619
rect -5976 610 -5716 616
rect -5660 616 -5654 619
rect -5406 616 -5400 619
rect -5660 610 -5400 616
rect -5344 616 -5338 619
rect -5090 616 -5084 619
rect -5344 610 -5084 616
rect -5028 616 -5022 619
rect -4774 616 -4768 619
rect -5028 610 -4768 616
rect -4712 616 -4706 619
rect -4458 616 -4452 619
rect -4712 610 -4452 616
rect -4396 616 -4390 619
rect -4142 616 -4136 619
rect -4396 610 -4136 616
rect -4080 616 -4074 619
rect -3826 616 -3820 619
rect -4080 610 -3820 616
rect -3764 616 -3758 619
rect -3510 616 -3504 619
rect -3764 610 -3504 616
rect -3448 616 -3442 619
rect -3194 616 -3188 619
rect -3448 610 -3188 616
rect -3132 616 -3126 619
rect -2878 616 -2872 619
rect -3132 610 -2872 616
rect -2816 616 -2810 619
rect -2562 616 -2556 619
rect -2816 610 -2556 616
rect -2500 616 -2494 619
rect -2246 616 -2240 619
rect -2500 610 -2240 616
rect -2184 616 -2178 619
rect -1930 616 -1924 619
rect -2184 610 -1924 616
rect -1868 616 -1862 619
rect -1614 616 -1608 619
rect -1868 610 -1608 616
rect -1552 616 -1546 619
rect -1298 616 -1292 619
rect -1552 610 -1292 616
rect -1236 616 -1230 619
rect -982 616 -976 619
rect -1236 610 -976 616
rect -920 616 -914 619
rect -666 616 -660 619
rect -920 610 -660 616
rect -604 616 -598 619
rect -350 616 -344 619
rect -604 610 -344 616
rect -288 616 -282 619
rect -34 616 -28 619
rect -288 610 -28 616
rect 28 616 34 619
rect 282 616 288 619
rect 28 610 288 616
rect 344 616 350 619
rect 598 616 604 619
rect 344 610 604 616
rect 660 616 666 619
rect 914 616 920 619
rect 660 610 920 616
rect 976 616 982 619
rect 1230 616 1236 619
rect 976 610 1236 616
rect 1292 616 1298 619
rect 1546 616 1552 619
rect 1292 610 1552 616
rect 1608 616 1614 619
rect 1862 616 1868 619
rect 1608 610 1868 616
rect 1924 616 1930 619
rect 2178 616 2184 619
rect 1924 610 2184 616
rect 2240 616 2246 619
rect 2494 616 2500 619
rect 2240 610 2500 616
rect 2556 616 2562 619
rect 2810 616 2816 619
rect 2556 610 2816 616
rect 2872 616 2878 619
rect 3126 616 3132 619
rect 2872 610 3132 616
rect 3188 616 3194 619
rect 3442 616 3448 619
rect 3188 610 3448 616
rect 3504 616 3510 619
rect 3758 616 3764 619
rect 3504 610 3764 616
rect 3820 616 3826 619
rect 4074 616 4080 619
rect 3820 610 4080 616
rect 4136 616 4142 619
rect 4390 616 4396 619
rect 4136 610 4396 616
rect 4452 616 4458 619
rect 4706 616 4712 619
rect 4452 610 4712 616
rect 4768 616 4774 619
rect 5022 616 5028 619
rect 4768 610 5028 616
rect 5084 616 5090 619
rect 5338 616 5344 619
rect 5084 610 5344 616
rect 5400 616 5406 619
rect 5654 616 5660 619
rect 5400 610 5660 616
rect 5716 616 5722 619
rect 5970 616 5976 619
rect 5716 610 5976 616
rect 6032 616 6038 619
rect 6286 616 6292 619
rect 6032 610 6292 616
rect 6348 616 6354 619
rect 6602 616 6608 619
rect 6348 610 6608 616
rect 6664 616 6670 619
rect 6918 616 6924 619
rect 6664 610 6924 616
rect 6980 616 6986 619
rect 7234 616 7240 619
rect 6980 610 7240 616
rect 7296 616 7302 619
rect 7550 616 7556 619
rect 7296 610 7556 616
rect 7612 616 7618 619
rect 7866 616 7872 619
rect 7612 610 7872 616
rect 7928 616 7934 619
rect 8182 616 8188 619
rect 7928 610 8188 616
rect 8244 616 8250 619
rect 8498 616 8504 619
rect 8244 610 8504 616
rect 8560 616 8566 619
rect 8814 616 8820 619
rect 8560 610 8820 616
rect 8876 616 8882 619
rect 9130 616 9136 619
rect 8876 610 9136 616
rect 9192 616 9198 619
rect 9446 616 9452 619
rect 9192 610 9452 616
rect 9508 616 9514 619
rect 9762 616 9768 619
rect 9508 610 9768 616
rect 9824 616 9830 619
rect 10078 616 10084 619
rect 9824 610 10084 616
rect 10140 616 10146 619
rect 10394 616 10400 619
rect 10140 610 10400 616
rect 10456 616 10462 619
rect 10710 616 10716 619
rect 10456 610 10716 616
rect 10772 616 10778 619
rect 11026 616 11032 619
rect 10772 610 11032 616
rect 11088 616 11094 619
rect 11342 616 11348 619
rect 11088 610 11348 616
rect 11404 616 11410 619
rect 11658 616 11664 619
rect 11404 610 11664 616
rect 11720 616 11726 619
rect 11974 616 11980 619
rect 11720 610 11980 616
rect 12036 616 12042 619
rect 12290 616 12296 619
rect 12036 610 12296 616
rect 12352 616 12358 619
rect 12606 616 12612 619
rect 12352 610 12612 616
rect 12668 616 12674 619
rect 12922 616 12928 619
rect 12668 610 12928 616
rect 12984 616 12990 619
rect 12984 610 13119 616
rect -13119 576 -13107 610
rect 13107 576 13119 610
rect -13119 570 -12984 576
rect -12990 567 -12984 570
rect -12928 570 -12668 576
rect -12928 567 -12922 570
rect -12674 567 -12668 570
rect -12612 570 -12352 576
rect -12612 567 -12606 570
rect -12358 567 -12352 570
rect -12296 570 -12036 576
rect -12296 567 -12290 570
rect -12042 567 -12036 570
rect -11980 570 -11720 576
rect -11980 567 -11974 570
rect -11726 567 -11720 570
rect -11664 570 -11404 576
rect -11664 567 -11658 570
rect -11410 567 -11404 570
rect -11348 570 -11088 576
rect -11348 567 -11342 570
rect -11094 567 -11088 570
rect -11032 570 -10772 576
rect -11032 567 -11026 570
rect -10778 567 -10772 570
rect -10716 570 -10456 576
rect -10716 567 -10710 570
rect -10462 567 -10456 570
rect -10400 570 -10140 576
rect -10400 567 -10394 570
rect -10146 567 -10140 570
rect -10084 570 -9824 576
rect -10084 567 -10078 570
rect -9830 567 -9824 570
rect -9768 570 -9508 576
rect -9768 567 -9762 570
rect -9514 567 -9508 570
rect -9452 570 -9192 576
rect -9452 567 -9446 570
rect -9198 567 -9192 570
rect -9136 570 -8876 576
rect -9136 567 -9130 570
rect -8882 567 -8876 570
rect -8820 570 -8560 576
rect -8820 567 -8814 570
rect -8566 567 -8560 570
rect -8504 570 -8244 576
rect -8504 567 -8498 570
rect -8250 567 -8244 570
rect -8188 570 -7928 576
rect -8188 567 -8182 570
rect -7934 567 -7928 570
rect -7872 570 -7612 576
rect -7872 567 -7866 570
rect -7618 567 -7612 570
rect -7556 570 -7296 576
rect -7556 567 -7550 570
rect -7302 567 -7296 570
rect -7240 570 -6980 576
rect -7240 567 -7234 570
rect -6986 567 -6980 570
rect -6924 570 -6664 576
rect -6924 567 -6918 570
rect -6670 567 -6664 570
rect -6608 570 -6348 576
rect -6608 567 -6602 570
rect -6354 567 -6348 570
rect -6292 570 -6032 576
rect -6292 567 -6286 570
rect -6038 567 -6032 570
rect -5976 570 -5716 576
rect -5976 567 -5970 570
rect -5722 567 -5716 570
rect -5660 570 -5400 576
rect -5660 567 -5654 570
rect -5406 567 -5400 570
rect -5344 570 -5084 576
rect -5344 567 -5338 570
rect -5090 567 -5084 570
rect -5028 570 -4768 576
rect -5028 567 -5022 570
rect -4774 567 -4768 570
rect -4712 570 -4452 576
rect -4712 567 -4706 570
rect -4458 567 -4452 570
rect -4396 570 -4136 576
rect -4396 567 -4390 570
rect -4142 567 -4136 570
rect -4080 570 -3820 576
rect -4080 567 -4074 570
rect -3826 567 -3820 570
rect -3764 570 -3504 576
rect -3764 567 -3758 570
rect -3510 567 -3504 570
rect -3448 570 -3188 576
rect -3448 567 -3442 570
rect -3194 567 -3188 570
rect -3132 570 -2872 576
rect -3132 567 -3126 570
rect -2878 567 -2872 570
rect -2816 570 -2556 576
rect -2816 567 -2810 570
rect -2562 567 -2556 570
rect -2500 570 -2240 576
rect -2500 567 -2494 570
rect -2246 567 -2240 570
rect -2184 570 -1924 576
rect -2184 567 -2178 570
rect -1930 567 -1924 570
rect -1868 570 -1608 576
rect -1868 567 -1862 570
rect -1614 567 -1608 570
rect -1552 570 -1292 576
rect -1552 567 -1546 570
rect -1298 567 -1292 570
rect -1236 570 -976 576
rect -1236 567 -1230 570
rect -982 567 -976 570
rect -920 570 -660 576
rect -920 567 -914 570
rect -666 567 -660 570
rect -604 570 -344 576
rect -604 567 -598 570
rect -350 567 -344 570
rect -288 570 -28 576
rect -288 567 -282 570
rect -34 567 -28 570
rect 28 570 288 576
rect 28 567 34 570
rect 282 567 288 570
rect 344 570 604 576
rect 344 567 350 570
rect 598 567 604 570
rect 660 570 920 576
rect 660 567 666 570
rect 914 567 920 570
rect 976 570 1236 576
rect 976 567 982 570
rect 1230 567 1236 570
rect 1292 570 1552 576
rect 1292 567 1298 570
rect 1546 567 1552 570
rect 1608 570 1868 576
rect 1608 567 1614 570
rect 1862 567 1868 570
rect 1924 570 2184 576
rect 1924 567 1930 570
rect 2178 567 2184 570
rect 2240 570 2500 576
rect 2240 567 2246 570
rect 2494 567 2500 570
rect 2556 570 2816 576
rect 2556 567 2562 570
rect 2810 567 2816 570
rect 2872 570 3132 576
rect 2872 567 2878 570
rect 3126 567 3132 570
rect 3188 570 3448 576
rect 3188 567 3194 570
rect 3442 567 3448 570
rect 3504 570 3764 576
rect 3504 567 3510 570
rect 3758 567 3764 570
rect 3820 570 4080 576
rect 3820 567 3826 570
rect 4074 567 4080 570
rect 4136 570 4396 576
rect 4136 567 4142 570
rect 4390 567 4396 570
rect 4452 570 4712 576
rect 4452 567 4458 570
rect 4706 567 4712 570
rect 4768 570 5028 576
rect 4768 567 4774 570
rect 5022 567 5028 570
rect 5084 570 5344 576
rect 5084 567 5090 570
rect 5338 567 5344 570
rect 5400 570 5660 576
rect 5400 567 5406 570
rect 5654 567 5660 570
rect 5716 570 5976 576
rect 5716 567 5722 570
rect 5970 567 5976 570
rect 6032 570 6292 576
rect 6032 567 6038 570
rect 6286 567 6292 570
rect 6348 570 6608 576
rect 6348 567 6354 570
rect 6602 567 6608 570
rect 6664 570 6924 576
rect 6664 567 6670 570
rect 6918 567 6924 570
rect 6980 570 7240 576
rect 6980 567 6986 570
rect 7234 567 7240 570
rect 7296 570 7556 576
rect 7296 567 7302 570
rect 7550 567 7556 570
rect 7612 570 7872 576
rect 7612 567 7618 570
rect 7866 567 7872 570
rect 7928 570 8188 576
rect 7928 567 7934 570
rect 8182 567 8188 570
rect 8244 570 8504 576
rect 8244 567 8250 570
rect 8498 567 8504 570
rect 8560 570 8820 576
rect 8560 567 8566 570
rect 8814 567 8820 570
rect 8876 570 9136 576
rect 8876 567 8882 570
rect 9130 567 9136 570
rect 9192 570 9452 576
rect 9192 567 9198 570
rect 9446 567 9452 570
rect 9508 570 9768 576
rect 9508 567 9514 570
rect 9762 567 9768 570
rect 9824 570 10084 576
rect 9824 567 9830 570
rect 10078 567 10084 570
rect 10140 570 10400 576
rect 10140 567 10146 570
rect 10394 567 10400 570
rect 10456 570 10716 576
rect 10456 567 10462 570
rect 10710 567 10716 570
rect 10772 570 11032 576
rect 10772 567 10778 570
rect 11026 567 11032 570
rect 11088 570 11348 576
rect 11088 567 11094 570
rect 11342 567 11348 570
rect 11404 570 11664 576
rect 11404 567 11410 570
rect 11658 567 11664 570
rect 11720 570 11980 576
rect 11720 567 11726 570
rect 11974 567 11980 570
rect 12036 570 12296 576
rect 12036 567 12042 570
rect 12290 567 12296 570
rect 12352 570 12612 576
rect 12352 567 12358 570
rect 12606 567 12612 570
rect 12668 570 12928 576
rect 12668 567 12674 570
rect 12922 567 12928 570
rect 12984 570 13119 576
rect 12984 567 12990 570
rect -13120 472 13120 524
rect -13120 438 -12911 472
rect -12843 438 -12753 472
rect -12685 438 -12595 472
rect -12527 438 -12437 472
rect -12369 438 -12279 472
rect -12211 438 -12121 472
rect -12053 438 -11963 472
rect -11895 438 -11805 472
rect -11737 438 -11647 472
rect -11579 438 -11489 472
rect -11421 438 -11331 472
rect -11263 438 -11173 472
rect -11105 438 -11015 472
rect -10947 438 -10857 472
rect -10789 438 -10699 472
rect -10631 438 -10541 472
rect -10473 438 -10383 472
rect -10315 438 -10225 472
rect -10157 438 -10067 472
rect -9999 438 -9909 472
rect -9841 438 -9751 472
rect -9683 438 -9593 472
rect -9525 438 -9435 472
rect -9367 438 -9277 472
rect -9209 438 -9119 472
rect -9051 438 -8961 472
rect -8893 438 -8803 472
rect -8735 438 -8645 472
rect -8577 438 -8487 472
rect -8419 438 -8329 472
rect -8261 438 -8171 472
rect -8103 438 -8013 472
rect -7945 438 -7855 472
rect -7787 438 -7697 472
rect -7629 438 -7539 472
rect -7471 438 -7381 472
rect -7313 438 -7223 472
rect -7155 438 -7065 472
rect -6997 438 -6907 472
rect -6839 438 -6749 472
rect -6681 438 -6591 472
rect -6523 438 -6433 472
rect -6365 438 -6275 472
rect -6207 438 -6117 472
rect -6049 438 -5959 472
rect -5891 438 -5801 472
rect -5733 438 -5643 472
rect -5575 438 -5485 472
rect -5417 438 -5327 472
rect -5259 438 -5169 472
rect -5101 438 -5011 472
rect -4943 438 -4853 472
rect -4785 438 -4695 472
rect -4627 438 -4537 472
rect -4469 438 -4379 472
rect -4311 438 -4221 472
rect -4153 438 -4063 472
rect -3995 438 -3905 472
rect -3837 438 -3747 472
rect -3679 438 -3589 472
rect -3521 438 -3431 472
rect -3363 438 -3273 472
rect -3205 438 -3115 472
rect -3047 438 -2957 472
rect -2889 438 -2799 472
rect -2731 438 -2641 472
rect -2573 438 -2483 472
rect -2415 438 -2325 472
rect -2257 438 -2167 472
rect -2099 438 -2009 472
rect -1941 438 -1851 472
rect -1783 438 -1693 472
rect -1625 438 -1535 472
rect -1467 438 -1377 472
rect -1309 438 -1219 472
rect -1151 438 -1061 472
rect -993 438 -903 472
rect -835 438 -745 472
rect -677 438 -587 472
rect -519 438 -429 472
rect -361 438 -271 472
rect -203 438 -113 472
rect -45 438 45 472
rect 113 438 203 472
rect 271 438 361 472
rect 429 438 519 472
rect 587 438 677 472
rect 745 438 835 472
rect 903 438 993 472
rect 1061 438 1151 472
rect 1219 438 1309 472
rect 1377 438 1467 472
rect 1535 438 1625 472
rect 1693 438 1783 472
rect 1851 438 1941 472
rect 2009 438 2099 472
rect 2167 438 2257 472
rect 2325 438 2415 472
rect 2483 438 2573 472
rect 2641 438 2731 472
rect 2799 438 2889 472
rect 2957 438 3047 472
rect 3115 438 3205 472
rect 3273 438 3363 472
rect 3431 438 3521 472
rect 3589 438 3679 472
rect 3747 438 3837 472
rect 3905 438 3995 472
rect 4063 438 4153 472
rect 4221 438 4311 472
rect 4379 438 4469 472
rect 4537 438 4627 472
rect 4695 438 4785 472
rect 4853 438 4943 472
rect 5011 438 5101 472
rect 5169 438 5259 472
rect 5327 438 5417 472
rect 5485 438 5575 472
rect 5643 438 5733 472
rect 5801 438 5891 472
rect 5959 438 6049 472
rect 6117 438 6207 472
rect 6275 438 6365 472
rect 6433 438 6523 472
rect 6591 438 6681 472
rect 6749 438 6839 472
rect 6907 438 6997 472
rect 7065 438 7155 472
rect 7223 438 7313 472
rect 7381 438 7471 472
rect 7539 438 7629 472
rect 7697 438 7787 472
rect 7855 438 7945 472
rect 8013 438 8103 472
rect 8171 438 8261 472
rect 8329 438 8419 472
rect 8487 438 8577 472
rect 8645 438 8735 472
rect 8803 438 8893 472
rect 8961 438 9051 472
rect 9119 438 9209 472
rect 9277 438 9367 472
rect 9435 438 9525 472
rect 9593 438 9683 472
rect 9751 438 9841 472
rect 9909 438 9999 472
rect 10067 438 10157 472
rect 10225 438 10315 472
rect 10383 438 10473 472
rect 10541 438 10631 472
rect 10699 438 10789 472
rect 10857 438 10947 472
rect 11015 438 11105 472
rect 11173 438 11263 472
rect 11331 438 11421 472
rect 11489 438 11579 472
rect 11647 438 11737 472
rect 11805 438 11895 472
rect 11963 438 12053 472
rect 12121 438 12211 472
rect 12279 438 12369 472
rect 12437 438 12527 472
rect 12595 438 12685 472
rect 12753 438 12843 472
rect 12911 438 13120 472
rect -13120 432 13120 438
rect -13120 -432 -13028 432
rect -12982 394 -12930 400
rect -12982 -400 -12930 -394
rect -12824 394 -12772 400
rect -12824 -400 -12772 -394
rect -12666 394 -12614 400
rect -12666 -400 -12614 -394
rect -12508 394 -12456 400
rect -12508 -400 -12456 -394
rect -12350 394 -12298 400
rect -12350 -400 -12298 -394
rect -12192 394 -12140 400
rect -12192 -400 -12140 -394
rect -12034 394 -11982 400
rect -12034 -400 -11982 -394
rect -11876 394 -11824 400
rect -11876 -400 -11824 -394
rect -11718 394 -11666 400
rect -11718 -400 -11666 -394
rect -11560 394 -11508 400
rect -11560 -400 -11508 -394
rect -11402 394 -11350 400
rect -11402 -400 -11350 -394
rect -11244 394 -11192 400
rect -11244 -400 -11192 -394
rect -11086 394 -11034 400
rect -11086 -400 -11034 -394
rect -10928 394 -10876 400
rect -10928 -400 -10876 -394
rect -10770 394 -10718 400
rect -10770 -400 -10718 -394
rect -10612 394 -10560 400
rect -10612 -400 -10560 -394
rect -10454 394 -10402 400
rect -10454 -400 -10402 -394
rect -10296 394 -10244 400
rect -10296 -400 -10244 -394
rect -10138 394 -10086 400
rect -10138 -400 -10086 -394
rect -9980 394 -9928 400
rect -9980 -400 -9928 -394
rect -9822 394 -9770 400
rect -9822 -400 -9770 -394
rect -9664 394 -9612 400
rect -9664 -400 -9612 -394
rect -9506 394 -9454 400
rect -9506 -400 -9454 -394
rect -9348 394 -9296 400
rect -9348 -400 -9296 -394
rect -9190 394 -9138 400
rect -9190 -400 -9138 -394
rect -9032 394 -8980 400
rect -9032 -400 -8980 -394
rect -8874 394 -8822 400
rect -8874 -400 -8822 -394
rect -8716 394 -8664 400
rect -8716 -400 -8664 -394
rect -8558 394 -8506 400
rect -8558 -400 -8506 -394
rect -8400 394 -8348 400
rect -8400 -400 -8348 -394
rect -8242 394 -8190 400
rect -8242 -400 -8190 -394
rect -8084 394 -8032 400
rect -8084 -400 -8032 -394
rect -7926 394 -7874 400
rect -7926 -400 -7874 -394
rect -7768 394 -7716 400
rect -7768 -400 -7716 -394
rect -7610 394 -7558 400
rect -7610 -400 -7558 -394
rect -7452 394 -7400 400
rect -7452 -400 -7400 -394
rect -7294 394 -7242 400
rect -7294 -400 -7242 -394
rect -7136 394 -7084 400
rect -7136 -400 -7084 -394
rect -6978 394 -6926 400
rect -6978 -400 -6926 -394
rect -6820 394 -6768 400
rect -6820 -400 -6768 -394
rect -6662 394 -6610 400
rect -6662 -400 -6610 -394
rect -6504 394 -6452 400
rect -6504 -400 -6452 -394
rect -6346 394 -6294 400
rect -6346 -400 -6294 -394
rect -6188 394 -6136 400
rect -6188 -400 -6136 -394
rect -6030 394 -5978 400
rect -6030 -400 -5978 -394
rect -5872 394 -5820 400
rect -5872 -400 -5820 -394
rect -5714 394 -5662 400
rect -5714 -400 -5662 -394
rect -5556 394 -5504 400
rect -5556 -400 -5504 -394
rect -5398 394 -5346 400
rect -5398 -400 -5346 -394
rect -5240 394 -5188 400
rect -5240 -400 -5188 -394
rect -5082 394 -5030 400
rect -5082 -400 -5030 -394
rect -4924 394 -4872 400
rect -4924 -400 -4872 -394
rect -4766 394 -4714 400
rect -4766 -400 -4714 -394
rect -4608 388 -4556 432
rect -4608 -388 -4599 388
rect -4565 -388 -4556 388
rect -4608 -432 -4556 -388
rect -4450 394 -4398 400
rect -4450 -400 -4398 -394
rect -4292 394 -4240 400
rect -4292 -400 -4240 -394
rect -4134 394 -4082 400
rect -4134 -400 -4082 -394
rect -3976 394 -3924 400
rect -3976 -400 -3924 -394
rect -3818 394 -3766 400
rect -3818 -400 -3766 -394
rect -3660 394 -3608 400
rect -3660 -400 -3608 -394
rect -3502 394 -3450 400
rect -3502 -400 -3450 -394
rect -3344 394 -3292 400
rect -3344 -400 -3292 -394
rect -3186 394 -3134 400
rect -3186 -400 -3134 -394
rect -3028 394 -2976 400
rect -3028 -400 -2976 -394
rect -2870 394 -2818 400
rect -2870 -400 -2818 -394
rect -2712 394 -2660 400
rect -2712 -400 -2660 -394
rect -2554 394 -2502 400
rect -2554 -400 -2502 -394
rect -2396 394 -2344 400
rect -2396 -400 -2344 -394
rect -2238 394 -2186 400
rect -2238 -400 -2186 -394
rect -2080 394 -2028 400
rect -2080 -400 -2028 -394
rect -1922 394 -1870 400
rect -1922 -400 -1870 -394
rect -1764 394 -1712 400
rect -1764 -400 -1712 -394
rect -1606 394 -1554 400
rect -1606 -400 -1554 -394
rect -1448 394 -1396 400
rect -1448 -400 -1396 -394
rect -1290 394 -1238 400
rect -1290 -400 -1238 -394
rect -1132 394 -1080 400
rect -1132 -400 -1080 -394
rect -974 394 -922 400
rect -974 -400 -922 -394
rect -816 394 -764 400
rect -816 -400 -764 -394
rect -658 394 -606 400
rect -658 -400 -606 -394
rect -500 394 -448 400
rect -500 -400 -448 -394
rect -342 394 -290 400
rect -342 -400 -290 -394
rect -184 394 -132 400
rect -184 -400 -132 -394
rect -26 394 26 400
rect -26 -400 26 -394
rect 132 394 184 400
rect 132 -400 184 -394
rect 290 394 342 400
rect 290 -400 342 -394
rect 448 394 500 400
rect 448 -400 500 -394
rect 606 394 658 400
rect 606 -400 658 -394
rect 764 394 816 400
rect 764 -400 816 -394
rect 922 394 974 400
rect 922 -400 974 -394
rect 1080 394 1132 400
rect 1080 -400 1132 -394
rect 1238 394 1290 400
rect 1238 -400 1290 -394
rect 1396 394 1448 400
rect 1396 -400 1448 -394
rect 1554 394 1606 400
rect 1554 -400 1606 -394
rect 1712 394 1764 400
rect 1712 -400 1764 -394
rect 1870 394 1922 400
rect 1870 -400 1922 -394
rect 2028 394 2080 400
rect 2028 -400 2080 -394
rect 2186 394 2238 400
rect 2186 -400 2238 -394
rect 2344 394 2396 400
rect 2344 -400 2396 -394
rect 2502 394 2554 400
rect 2502 -400 2554 -394
rect 2660 394 2712 400
rect 2660 -400 2712 -394
rect 2818 394 2870 400
rect 2818 -400 2870 -394
rect 2976 394 3028 400
rect 2976 -400 3028 -394
rect 3134 394 3186 400
rect 3134 -400 3186 -394
rect 3292 394 3344 400
rect 3292 -400 3344 -394
rect 3450 394 3502 400
rect 3450 -400 3502 -394
rect 3608 394 3660 400
rect 3608 -400 3660 -394
rect 3766 394 3818 400
rect 3766 -400 3818 -394
rect 3924 394 3976 400
rect 3924 -400 3976 -394
rect 4082 394 4134 400
rect 4082 -400 4134 -394
rect 4240 394 4292 400
rect 4240 -400 4292 -394
rect 4398 394 4450 400
rect 4398 -400 4450 -394
rect 4556 388 4608 432
rect 4556 -388 4565 388
rect 4599 -388 4608 388
rect 4556 -432 4608 -388
rect 4714 394 4766 400
rect 4714 -400 4766 -394
rect 4872 394 4924 400
rect 4872 -400 4924 -394
rect 5030 394 5082 400
rect 5030 -400 5082 -394
rect 5188 394 5240 400
rect 5188 -400 5240 -394
rect 5346 394 5398 400
rect 5346 -400 5398 -394
rect 5504 394 5556 400
rect 5504 -400 5556 -394
rect 5662 394 5714 400
rect 5662 -400 5714 -394
rect 5820 394 5872 400
rect 5820 -400 5872 -394
rect 5978 394 6030 400
rect 5978 -400 6030 -394
rect 6136 394 6188 400
rect 6136 -400 6188 -394
rect 6294 394 6346 400
rect 6294 -400 6346 -394
rect 6452 394 6504 400
rect 6452 -400 6504 -394
rect 6610 394 6662 400
rect 6610 -400 6662 -394
rect 6768 394 6820 400
rect 6768 -400 6820 -394
rect 6926 394 6978 400
rect 6926 -400 6978 -394
rect 7084 394 7136 400
rect 7084 -400 7136 -394
rect 7242 394 7294 400
rect 7242 -400 7294 -394
rect 7400 394 7452 400
rect 7400 -400 7452 -394
rect 7558 394 7610 400
rect 7558 -400 7610 -394
rect 7716 394 7768 400
rect 7716 -400 7768 -394
rect 7874 394 7926 400
rect 7874 -400 7926 -394
rect 8032 394 8084 400
rect 8032 -400 8084 -394
rect 8190 394 8242 400
rect 8190 -400 8242 -394
rect 8348 394 8400 400
rect 8348 -400 8400 -394
rect 8506 394 8558 400
rect 8506 -400 8558 -394
rect 8664 394 8716 400
rect 8664 -400 8716 -394
rect 8822 394 8874 400
rect 8822 -400 8874 -394
rect 8980 394 9032 400
rect 8980 -400 9032 -394
rect 9138 394 9190 400
rect 9138 -400 9190 -394
rect 9296 394 9348 400
rect 9296 -400 9348 -394
rect 9454 394 9506 400
rect 9454 -400 9506 -394
rect 9612 394 9664 400
rect 9612 -400 9664 -394
rect 9770 394 9822 400
rect 9770 -400 9822 -394
rect 9928 394 9980 400
rect 9928 -400 9980 -394
rect 10086 394 10138 400
rect 10086 -400 10138 -394
rect 10244 394 10296 400
rect 10244 -400 10296 -394
rect 10402 394 10454 400
rect 10402 -400 10454 -394
rect 10560 394 10612 400
rect 10560 -400 10612 -394
rect 10718 394 10770 400
rect 10718 -400 10770 -394
rect 10876 394 10928 400
rect 10876 -400 10928 -394
rect 11034 394 11086 400
rect 11034 -400 11086 -394
rect 11192 394 11244 400
rect 11192 -400 11244 -394
rect 11350 394 11402 400
rect 11350 -400 11402 -394
rect 11508 394 11560 400
rect 11508 -400 11560 -394
rect 11666 394 11718 400
rect 11666 -400 11718 -394
rect 11824 394 11876 400
rect 11824 -400 11876 -394
rect 11982 394 12034 400
rect 11982 -400 12034 -394
rect 12140 394 12192 400
rect 12140 -400 12192 -394
rect 12298 394 12350 400
rect 12298 -400 12350 -394
rect 12456 394 12508 400
rect 12456 -400 12508 -394
rect 12614 394 12666 400
rect 12614 -400 12666 -394
rect 12772 394 12824 400
rect 12772 -400 12824 -394
rect 12930 394 12982 400
rect 12930 -400 12982 -394
rect 13028 -432 13120 432
rect -13120 -438 13120 -432
rect -13120 -472 -12911 -438
rect -12843 -472 -12753 -438
rect -12685 -472 -12595 -438
rect -12527 -472 -12437 -438
rect -12369 -472 -12279 -438
rect -12211 -472 -12121 -438
rect -12053 -472 -11963 -438
rect -11895 -472 -11805 -438
rect -11737 -472 -11647 -438
rect -11579 -472 -11489 -438
rect -11421 -472 -11331 -438
rect -11263 -472 -11173 -438
rect -11105 -472 -11015 -438
rect -10947 -472 -10857 -438
rect -10789 -472 -10699 -438
rect -10631 -472 -10541 -438
rect -10473 -472 -10383 -438
rect -10315 -472 -10225 -438
rect -10157 -472 -10067 -438
rect -9999 -472 -9909 -438
rect -9841 -472 -9751 -438
rect -9683 -472 -9593 -438
rect -9525 -472 -9435 -438
rect -9367 -472 -9277 -438
rect -9209 -472 -9119 -438
rect -9051 -472 -8961 -438
rect -8893 -472 -8803 -438
rect -8735 -472 -8645 -438
rect -8577 -472 -8487 -438
rect -8419 -472 -8329 -438
rect -8261 -472 -8171 -438
rect -8103 -472 -8013 -438
rect -7945 -472 -7855 -438
rect -7787 -472 -7697 -438
rect -7629 -472 -7539 -438
rect -7471 -472 -7381 -438
rect -7313 -472 -7223 -438
rect -7155 -472 -7065 -438
rect -6997 -472 -6907 -438
rect -6839 -472 -6749 -438
rect -6681 -472 -6591 -438
rect -6523 -472 -6433 -438
rect -6365 -472 -6275 -438
rect -6207 -472 -6117 -438
rect -6049 -472 -5959 -438
rect -5891 -472 -5801 -438
rect -5733 -472 -5643 -438
rect -5575 -472 -5485 -438
rect -5417 -472 -5327 -438
rect -5259 -472 -5169 -438
rect -5101 -472 -5011 -438
rect -4943 -472 -4853 -438
rect -4785 -472 -4695 -438
rect -4627 -472 -4537 -438
rect -4469 -472 -4379 -438
rect -4311 -472 -4221 -438
rect -4153 -472 -4063 -438
rect -3995 -472 -3905 -438
rect -3837 -472 -3747 -438
rect -3679 -472 -3589 -438
rect -3521 -472 -3431 -438
rect -3363 -472 -3273 -438
rect -3205 -472 -3115 -438
rect -3047 -472 -2957 -438
rect -2889 -472 -2799 -438
rect -2731 -472 -2641 -438
rect -2573 -472 -2483 -438
rect -2415 -472 -2325 -438
rect -2257 -472 -2167 -438
rect -2099 -472 -2009 -438
rect -1941 -472 -1851 -438
rect -1783 -472 -1693 -438
rect -1625 -472 -1535 -438
rect -1467 -472 -1377 -438
rect -1309 -472 -1219 -438
rect -1151 -472 -1061 -438
rect -993 -472 -903 -438
rect -835 -472 -745 -438
rect -677 -472 -587 -438
rect -519 -472 -429 -438
rect -361 -472 -271 -438
rect -203 -472 -113 -438
rect -45 -472 45 -438
rect 113 -472 203 -438
rect 271 -472 361 -438
rect 429 -472 519 -438
rect 587 -472 677 -438
rect 745 -472 835 -438
rect 903 -472 993 -438
rect 1061 -472 1151 -438
rect 1219 -472 1309 -438
rect 1377 -472 1467 -438
rect 1535 -472 1625 -438
rect 1693 -472 1783 -438
rect 1851 -472 1941 -438
rect 2009 -472 2099 -438
rect 2167 -472 2257 -438
rect 2325 -472 2415 -438
rect 2483 -472 2573 -438
rect 2641 -472 2731 -438
rect 2799 -472 2889 -438
rect 2957 -472 3047 -438
rect 3115 -472 3205 -438
rect 3273 -472 3363 -438
rect 3431 -472 3521 -438
rect 3589 -472 3679 -438
rect 3747 -472 3837 -438
rect 3905 -472 3995 -438
rect 4063 -472 4153 -438
rect 4221 -472 4311 -438
rect 4379 -472 4469 -438
rect 4537 -472 4627 -438
rect 4695 -472 4785 -438
rect 4853 -472 4943 -438
rect 5011 -472 5101 -438
rect 5169 -472 5259 -438
rect 5327 -472 5417 -438
rect 5485 -472 5575 -438
rect 5643 -472 5733 -438
rect 5801 -472 5891 -438
rect 5959 -472 6049 -438
rect 6117 -472 6207 -438
rect 6275 -472 6365 -438
rect 6433 -472 6523 -438
rect 6591 -472 6681 -438
rect 6749 -472 6839 -438
rect 6907 -472 6997 -438
rect 7065 -472 7155 -438
rect 7223 -472 7313 -438
rect 7381 -472 7471 -438
rect 7539 -472 7629 -438
rect 7697 -472 7787 -438
rect 7855 -472 7945 -438
rect 8013 -472 8103 -438
rect 8171 -472 8261 -438
rect 8329 -472 8419 -438
rect 8487 -472 8577 -438
rect 8645 -472 8735 -438
rect 8803 -472 8893 -438
rect 8961 -472 9051 -438
rect 9119 -472 9209 -438
rect 9277 -472 9367 -438
rect 9435 -472 9525 -438
rect 9593 -472 9683 -438
rect 9751 -472 9841 -438
rect 9909 -472 9999 -438
rect 10067 -472 10157 -438
rect 10225 -472 10315 -438
rect 10383 -472 10473 -438
rect 10541 -472 10631 -438
rect 10699 -472 10789 -438
rect 10857 -472 10947 -438
rect 11015 -472 11105 -438
rect 11173 -472 11263 -438
rect 11331 -472 11421 -438
rect 11489 -472 11579 -438
rect 11647 -472 11737 -438
rect 11805 -472 11895 -438
rect 11963 -472 12053 -438
rect 12121 -472 12211 -438
rect 12279 -472 12369 -438
rect 12437 -472 12527 -438
rect 12595 -472 12685 -438
rect 12753 -472 12843 -438
rect 12911 -472 13120 -438
rect -13120 -524 13120 -472
rect -12990 -570 -12984 -567
rect -13119 -576 -12984 -570
rect -12928 -570 -12922 -567
rect -12674 -570 -12668 -567
rect -12928 -576 -12668 -570
rect -12612 -570 -12606 -567
rect -12358 -570 -12352 -567
rect -12612 -576 -12352 -570
rect -12296 -570 -12290 -567
rect -12042 -570 -12036 -567
rect -12296 -576 -12036 -570
rect -11980 -570 -11974 -567
rect -11726 -570 -11720 -567
rect -11980 -576 -11720 -570
rect -11664 -570 -11658 -567
rect -11410 -570 -11404 -567
rect -11664 -576 -11404 -570
rect -11348 -570 -11342 -567
rect -11094 -570 -11088 -567
rect -11348 -576 -11088 -570
rect -11032 -570 -11026 -567
rect -10778 -570 -10772 -567
rect -11032 -576 -10772 -570
rect -10716 -570 -10710 -567
rect -10462 -570 -10456 -567
rect -10716 -576 -10456 -570
rect -10400 -570 -10394 -567
rect -10146 -570 -10140 -567
rect -10400 -576 -10140 -570
rect -10084 -570 -10078 -567
rect -9830 -570 -9824 -567
rect -10084 -576 -9824 -570
rect -9768 -570 -9762 -567
rect -9514 -570 -9508 -567
rect -9768 -576 -9508 -570
rect -9452 -570 -9446 -567
rect -9198 -570 -9192 -567
rect -9452 -576 -9192 -570
rect -9136 -570 -9130 -567
rect -8882 -570 -8876 -567
rect -9136 -576 -8876 -570
rect -8820 -570 -8814 -567
rect -8566 -570 -8560 -567
rect -8820 -576 -8560 -570
rect -8504 -570 -8498 -567
rect -8250 -570 -8244 -567
rect -8504 -576 -8244 -570
rect -8188 -570 -8182 -567
rect -7934 -570 -7928 -567
rect -8188 -576 -7928 -570
rect -7872 -570 -7866 -567
rect -7618 -570 -7612 -567
rect -7872 -576 -7612 -570
rect -7556 -570 -7550 -567
rect -7302 -570 -7296 -567
rect -7556 -576 -7296 -570
rect -7240 -570 -7234 -567
rect -6986 -570 -6980 -567
rect -7240 -576 -6980 -570
rect -6924 -570 -6918 -567
rect -6670 -570 -6664 -567
rect -6924 -576 -6664 -570
rect -6608 -570 -6602 -567
rect -6354 -570 -6348 -567
rect -6608 -576 -6348 -570
rect -6292 -570 -6286 -567
rect -6038 -570 -6032 -567
rect -6292 -576 -6032 -570
rect -5976 -570 -5970 -567
rect -5722 -570 -5716 -567
rect -5976 -576 -5716 -570
rect -5660 -570 -5654 -567
rect -5406 -570 -5400 -567
rect -5660 -576 -5400 -570
rect -5344 -570 -5338 -567
rect -5090 -570 -5084 -567
rect -5344 -576 -5084 -570
rect -5028 -570 -5022 -567
rect -4774 -570 -4768 -567
rect -5028 -576 -4768 -570
rect -4712 -570 -4706 -567
rect -4458 -570 -4452 -567
rect -4712 -576 -4452 -570
rect -4396 -570 -4390 -567
rect -4142 -570 -4136 -567
rect -4396 -576 -4136 -570
rect -4080 -570 -4074 -567
rect -3826 -570 -3820 -567
rect -4080 -576 -3820 -570
rect -3764 -570 -3758 -567
rect -3510 -570 -3504 -567
rect -3764 -576 -3504 -570
rect -3448 -570 -3442 -567
rect -3194 -570 -3188 -567
rect -3448 -576 -3188 -570
rect -3132 -570 -3126 -567
rect -2878 -570 -2872 -567
rect -3132 -576 -2872 -570
rect -2816 -570 -2810 -567
rect -2562 -570 -2556 -567
rect -2816 -576 -2556 -570
rect -2500 -570 -2494 -567
rect -2246 -570 -2240 -567
rect -2500 -576 -2240 -570
rect -2184 -570 -2178 -567
rect -1930 -570 -1924 -567
rect -2184 -576 -1924 -570
rect -1868 -570 -1862 -567
rect -1614 -570 -1608 -567
rect -1868 -576 -1608 -570
rect -1552 -570 -1546 -567
rect -1298 -570 -1292 -567
rect -1552 -576 -1292 -570
rect -1236 -570 -1230 -567
rect -982 -570 -976 -567
rect -1236 -576 -976 -570
rect -920 -570 -914 -567
rect -666 -570 -660 -567
rect -920 -576 -660 -570
rect -604 -570 -598 -567
rect -350 -570 -344 -567
rect -604 -576 -344 -570
rect -288 -570 -282 -567
rect -34 -570 -28 -567
rect -288 -576 -28 -570
rect 28 -570 34 -567
rect 282 -570 288 -567
rect 28 -576 288 -570
rect 344 -570 350 -567
rect 598 -570 604 -567
rect 344 -576 604 -570
rect 660 -570 666 -567
rect 914 -570 920 -567
rect 660 -576 920 -570
rect 976 -570 982 -567
rect 1230 -570 1236 -567
rect 976 -576 1236 -570
rect 1292 -570 1298 -567
rect 1546 -570 1552 -567
rect 1292 -576 1552 -570
rect 1608 -570 1614 -567
rect 1862 -570 1868 -567
rect 1608 -576 1868 -570
rect 1924 -570 1930 -567
rect 2178 -570 2184 -567
rect 1924 -576 2184 -570
rect 2240 -570 2246 -567
rect 2494 -570 2500 -567
rect 2240 -576 2500 -570
rect 2556 -570 2562 -567
rect 2810 -570 2816 -567
rect 2556 -576 2816 -570
rect 2872 -570 2878 -567
rect 3126 -570 3132 -567
rect 2872 -576 3132 -570
rect 3188 -570 3194 -567
rect 3442 -570 3448 -567
rect 3188 -576 3448 -570
rect 3504 -570 3510 -567
rect 3758 -570 3764 -567
rect 3504 -576 3764 -570
rect 3820 -570 3826 -567
rect 4074 -570 4080 -567
rect 3820 -576 4080 -570
rect 4136 -570 4142 -567
rect 4390 -570 4396 -567
rect 4136 -576 4396 -570
rect 4452 -570 4458 -567
rect 4706 -570 4712 -567
rect 4452 -576 4712 -570
rect 4768 -570 4774 -567
rect 5022 -570 5028 -567
rect 4768 -576 5028 -570
rect 5084 -570 5090 -567
rect 5338 -570 5344 -567
rect 5084 -576 5344 -570
rect 5400 -570 5406 -567
rect 5654 -570 5660 -567
rect 5400 -576 5660 -570
rect 5716 -570 5722 -567
rect 5970 -570 5976 -567
rect 5716 -576 5976 -570
rect 6032 -570 6038 -567
rect 6286 -570 6292 -567
rect 6032 -576 6292 -570
rect 6348 -570 6354 -567
rect 6602 -570 6608 -567
rect 6348 -576 6608 -570
rect 6664 -570 6670 -567
rect 6918 -570 6924 -567
rect 6664 -576 6924 -570
rect 6980 -570 6986 -567
rect 7234 -570 7240 -567
rect 6980 -576 7240 -570
rect 7296 -570 7302 -567
rect 7550 -570 7556 -567
rect 7296 -576 7556 -570
rect 7612 -570 7618 -567
rect 7866 -570 7872 -567
rect 7612 -576 7872 -570
rect 7928 -570 7934 -567
rect 8182 -570 8188 -567
rect 7928 -576 8188 -570
rect 8244 -570 8250 -567
rect 8498 -570 8504 -567
rect 8244 -576 8504 -570
rect 8560 -570 8566 -567
rect 8814 -570 8820 -567
rect 8560 -576 8820 -570
rect 8876 -570 8882 -567
rect 9130 -570 9136 -567
rect 8876 -576 9136 -570
rect 9192 -570 9198 -567
rect 9446 -570 9452 -567
rect 9192 -576 9452 -570
rect 9508 -570 9514 -567
rect 9762 -570 9768 -567
rect 9508 -576 9768 -570
rect 9824 -570 9830 -567
rect 10078 -570 10084 -567
rect 9824 -576 10084 -570
rect 10140 -570 10146 -567
rect 10394 -570 10400 -567
rect 10140 -576 10400 -570
rect 10456 -570 10462 -567
rect 10710 -570 10716 -567
rect 10456 -576 10716 -570
rect 10772 -570 10778 -567
rect 11026 -570 11032 -567
rect 10772 -576 11032 -570
rect 11088 -570 11094 -567
rect 11342 -570 11348 -567
rect 11088 -576 11348 -570
rect 11404 -570 11410 -567
rect 11658 -570 11664 -567
rect 11404 -576 11664 -570
rect 11720 -570 11726 -567
rect 11974 -570 11980 -567
rect 11720 -576 11980 -570
rect 12036 -570 12042 -567
rect 12290 -570 12296 -567
rect 12036 -576 12296 -570
rect 12352 -570 12358 -567
rect 12606 -570 12612 -567
rect 12352 -576 12612 -570
rect 12668 -570 12674 -567
rect 12922 -570 12928 -567
rect 12668 -576 12928 -570
rect 12984 -570 12990 -567
rect 12984 -576 13119 -570
rect -13119 -610 -13107 -576
rect 13107 -610 13119 -576
rect -13119 -616 -12984 -610
rect -12990 -619 -12984 -616
rect -12928 -616 -12668 -610
rect -12928 -619 -12922 -616
rect -12674 -619 -12668 -616
rect -12612 -616 -12352 -610
rect -12612 -619 -12606 -616
rect -12358 -619 -12352 -616
rect -12296 -616 -12036 -610
rect -12296 -619 -12290 -616
rect -12042 -619 -12036 -616
rect -11980 -616 -11720 -610
rect -11980 -619 -11974 -616
rect -11726 -619 -11720 -616
rect -11664 -616 -11404 -610
rect -11664 -619 -11658 -616
rect -11410 -619 -11404 -616
rect -11348 -616 -11088 -610
rect -11348 -619 -11342 -616
rect -11094 -619 -11088 -616
rect -11032 -616 -10772 -610
rect -11032 -619 -11026 -616
rect -10778 -619 -10772 -616
rect -10716 -616 -10456 -610
rect -10716 -619 -10710 -616
rect -10462 -619 -10456 -616
rect -10400 -616 -10140 -610
rect -10400 -619 -10394 -616
rect -10146 -619 -10140 -616
rect -10084 -616 -9824 -610
rect -10084 -619 -10078 -616
rect -9830 -619 -9824 -616
rect -9768 -616 -9508 -610
rect -9768 -619 -9762 -616
rect -9514 -619 -9508 -616
rect -9452 -616 -9192 -610
rect -9452 -619 -9446 -616
rect -9198 -619 -9192 -616
rect -9136 -616 -8876 -610
rect -9136 -619 -9130 -616
rect -8882 -619 -8876 -616
rect -8820 -616 -8560 -610
rect -8820 -619 -8814 -616
rect -8566 -619 -8560 -616
rect -8504 -616 -8244 -610
rect -8504 -619 -8498 -616
rect -8250 -619 -8244 -616
rect -8188 -616 -7928 -610
rect -8188 -619 -8182 -616
rect -7934 -619 -7928 -616
rect -7872 -616 -7612 -610
rect -7872 -619 -7866 -616
rect -7618 -619 -7612 -616
rect -7556 -616 -7296 -610
rect -7556 -619 -7550 -616
rect -7302 -619 -7296 -616
rect -7240 -616 -6980 -610
rect -7240 -619 -7234 -616
rect -6986 -619 -6980 -616
rect -6924 -616 -6664 -610
rect -6924 -619 -6918 -616
rect -6670 -619 -6664 -616
rect -6608 -616 -6348 -610
rect -6608 -619 -6602 -616
rect -6354 -619 -6348 -616
rect -6292 -616 -6032 -610
rect -6292 -619 -6286 -616
rect -6038 -619 -6032 -616
rect -5976 -616 -5716 -610
rect -5976 -619 -5970 -616
rect -5722 -619 -5716 -616
rect -5660 -616 -5400 -610
rect -5660 -619 -5654 -616
rect -5406 -619 -5400 -616
rect -5344 -616 -5084 -610
rect -5344 -619 -5338 -616
rect -5090 -619 -5084 -616
rect -5028 -616 -4768 -610
rect -5028 -619 -5022 -616
rect -4774 -619 -4768 -616
rect -4712 -616 -4452 -610
rect -4712 -619 -4706 -616
rect -4458 -619 -4452 -616
rect -4396 -616 -4136 -610
rect -4396 -619 -4390 -616
rect -4142 -619 -4136 -616
rect -4080 -616 -3820 -610
rect -4080 -619 -4074 -616
rect -3826 -619 -3820 -616
rect -3764 -616 -3504 -610
rect -3764 -619 -3758 -616
rect -3510 -619 -3504 -616
rect -3448 -616 -3188 -610
rect -3448 -619 -3442 -616
rect -3194 -619 -3188 -616
rect -3132 -616 -2872 -610
rect -3132 -619 -3126 -616
rect -2878 -619 -2872 -616
rect -2816 -616 -2556 -610
rect -2816 -619 -2810 -616
rect -2562 -619 -2556 -616
rect -2500 -616 -2240 -610
rect -2500 -619 -2494 -616
rect -2246 -619 -2240 -616
rect -2184 -616 -1924 -610
rect -2184 -619 -2178 -616
rect -1930 -619 -1924 -616
rect -1868 -616 -1608 -610
rect -1868 -619 -1862 -616
rect -1614 -619 -1608 -616
rect -1552 -616 -1292 -610
rect -1552 -619 -1546 -616
rect -1298 -619 -1292 -616
rect -1236 -616 -976 -610
rect -1236 -619 -1230 -616
rect -982 -619 -976 -616
rect -920 -616 -660 -610
rect -920 -619 -914 -616
rect -666 -619 -660 -616
rect -604 -616 -344 -610
rect -604 -619 -598 -616
rect -350 -619 -344 -616
rect -288 -616 -28 -610
rect -288 -619 -282 -616
rect -34 -619 -28 -616
rect 28 -616 288 -610
rect 28 -619 34 -616
rect 282 -619 288 -616
rect 344 -616 604 -610
rect 344 -619 350 -616
rect 598 -619 604 -616
rect 660 -616 920 -610
rect 660 -619 666 -616
rect 914 -619 920 -616
rect 976 -616 1236 -610
rect 976 -619 982 -616
rect 1230 -619 1236 -616
rect 1292 -616 1552 -610
rect 1292 -619 1298 -616
rect 1546 -619 1552 -616
rect 1608 -616 1868 -610
rect 1608 -619 1614 -616
rect 1862 -619 1868 -616
rect 1924 -616 2184 -610
rect 1924 -619 1930 -616
rect 2178 -619 2184 -616
rect 2240 -616 2500 -610
rect 2240 -619 2246 -616
rect 2494 -619 2500 -616
rect 2556 -616 2816 -610
rect 2556 -619 2562 -616
rect 2810 -619 2816 -616
rect 2872 -616 3132 -610
rect 2872 -619 2878 -616
rect 3126 -619 3132 -616
rect 3188 -616 3448 -610
rect 3188 -619 3194 -616
rect 3442 -619 3448 -616
rect 3504 -616 3764 -610
rect 3504 -619 3510 -616
rect 3758 -619 3764 -616
rect 3820 -616 4080 -610
rect 3820 -619 3826 -616
rect 4074 -619 4080 -616
rect 4136 -616 4396 -610
rect 4136 -619 4142 -616
rect 4390 -619 4396 -616
rect 4452 -616 4712 -610
rect 4452 -619 4458 -616
rect 4706 -619 4712 -616
rect 4768 -616 5028 -610
rect 4768 -619 4774 -616
rect 5022 -619 5028 -616
rect 5084 -616 5344 -610
rect 5084 -619 5090 -616
rect 5338 -619 5344 -616
rect 5400 -616 5660 -610
rect 5400 -619 5406 -616
rect 5654 -619 5660 -616
rect 5716 -616 5976 -610
rect 5716 -619 5722 -616
rect 5970 -619 5976 -616
rect 6032 -616 6292 -610
rect 6032 -619 6038 -616
rect 6286 -619 6292 -616
rect 6348 -616 6608 -610
rect 6348 -619 6354 -616
rect 6602 -619 6608 -616
rect 6664 -616 6924 -610
rect 6664 -619 6670 -616
rect 6918 -619 6924 -616
rect 6980 -616 7240 -610
rect 6980 -619 6986 -616
rect 7234 -619 7240 -616
rect 7296 -616 7556 -610
rect 7296 -619 7302 -616
rect 7550 -619 7556 -616
rect 7612 -616 7872 -610
rect 7612 -619 7618 -616
rect 7866 -619 7872 -616
rect 7928 -616 8188 -610
rect 7928 -619 7934 -616
rect 8182 -619 8188 -616
rect 8244 -616 8504 -610
rect 8244 -619 8250 -616
rect 8498 -619 8504 -616
rect 8560 -616 8820 -610
rect 8560 -619 8566 -616
rect 8814 -619 8820 -616
rect 8876 -616 9136 -610
rect 8876 -619 8882 -616
rect 9130 -619 9136 -616
rect 9192 -616 9452 -610
rect 9192 -619 9198 -616
rect 9446 -619 9452 -616
rect 9508 -616 9768 -610
rect 9508 -619 9514 -616
rect 9762 -619 9768 -616
rect 9824 -616 10084 -610
rect 9824 -619 9830 -616
rect 10078 -619 10084 -616
rect 10140 -616 10400 -610
rect 10140 -619 10146 -616
rect 10394 -619 10400 -616
rect 10456 -616 10716 -610
rect 10456 -619 10462 -616
rect 10710 -619 10716 -616
rect 10772 -616 11032 -610
rect 10772 -619 10778 -616
rect 11026 -619 11032 -616
rect 11088 -616 11348 -610
rect 11088 -619 11094 -616
rect 11342 -619 11348 -616
rect 11404 -616 11664 -610
rect 11404 -619 11410 -616
rect 11658 -619 11664 -616
rect 11720 -616 11980 -610
rect 11720 -619 11726 -616
rect 11974 -619 11980 -616
rect 12036 -616 12296 -610
rect 12036 -619 12042 -616
rect 12290 -619 12296 -616
rect 12352 -616 12612 -610
rect 12352 -619 12358 -616
rect 12606 -619 12612 -616
rect 12668 -616 12928 -610
rect 12668 -619 12674 -616
rect 12922 -619 12928 -616
rect 12984 -616 13119 -610
rect 12984 -619 12990 -616
<< via1 >>
rect -12984 610 -12928 619
rect -12668 610 -12612 619
rect -12352 610 -12296 619
rect -12036 610 -11980 619
rect -11720 610 -11664 619
rect -11404 610 -11348 619
rect -11088 610 -11032 619
rect -10772 610 -10716 619
rect -10456 610 -10400 619
rect -10140 610 -10084 619
rect -9824 610 -9768 619
rect -9508 610 -9452 619
rect -9192 610 -9136 619
rect -8876 610 -8820 619
rect -8560 610 -8504 619
rect -8244 610 -8188 619
rect -7928 610 -7872 619
rect -7612 610 -7556 619
rect -7296 610 -7240 619
rect -6980 610 -6924 619
rect -6664 610 -6608 619
rect -6348 610 -6292 619
rect -6032 610 -5976 619
rect -5716 610 -5660 619
rect -5400 610 -5344 619
rect -5084 610 -5028 619
rect -4768 610 -4712 619
rect -4452 610 -4396 619
rect -4136 610 -4080 619
rect -3820 610 -3764 619
rect -3504 610 -3448 619
rect -3188 610 -3132 619
rect -2872 610 -2816 619
rect -2556 610 -2500 619
rect -2240 610 -2184 619
rect -1924 610 -1868 619
rect -1608 610 -1552 619
rect -1292 610 -1236 619
rect -976 610 -920 619
rect -660 610 -604 619
rect -344 610 -288 619
rect -28 610 28 619
rect 288 610 344 619
rect 604 610 660 619
rect 920 610 976 619
rect 1236 610 1292 619
rect 1552 610 1608 619
rect 1868 610 1924 619
rect 2184 610 2240 619
rect 2500 610 2556 619
rect 2816 610 2872 619
rect 3132 610 3188 619
rect 3448 610 3504 619
rect 3764 610 3820 619
rect 4080 610 4136 619
rect 4396 610 4452 619
rect 4712 610 4768 619
rect 5028 610 5084 619
rect 5344 610 5400 619
rect 5660 610 5716 619
rect 5976 610 6032 619
rect 6292 610 6348 619
rect 6608 610 6664 619
rect 6924 610 6980 619
rect 7240 610 7296 619
rect 7556 610 7612 619
rect 7872 610 7928 619
rect 8188 610 8244 619
rect 8504 610 8560 619
rect 8820 610 8876 619
rect 9136 610 9192 619
rect 9452 610 9508 619
rect 9768 610 9824 619
rect 10084 610 10140 619
rect 10400 610 10456 619
rect 10716 610 10772 619
rect 11032 610 11088 619
rect 11348 610 11404 619
rect 11664 610 11720 619
rect 11980 610 12036 619
rect 12296 610 12352 619
rect 12612 610 12668 619
rect 12928 610 12984 619
rect -12984 576 -12928 610
rect -12668 576 -12612 610
rect -12352 576 -12296 610
rect -12036 576 -11980 610
rect -11720 576 -11664 610
rect -11404 576 -11348 610
rect -11088 576 -11032 610
rect -10772 576 -10716 610
rect -10456 576 -10400 610
rect -10140 576 -10084 610
rect -9824 576 -9768 610
rect -9508 576 -9452 610
rect -9192 576 -9136 610
rect -8876 576 -8820 610
rect -8560 576 -8504 610
rect -8244 576 -8188 610
rect -7928 576 -7872 610
rect -7612 576 -7556 610
rect -7296 576 -7240 610
rect -6980 576 -6924 610
rect -6664 576 -6608 610
rect -6348 576 -6292 610
rect -6032 576 -5976 610
rect -5716 576 -5660 610
rect -5400 576 -5344 610
rect -5084 576 -5028 610
rect -4768 576 -4712 610
rect -4452 576 -4396 610
rect -4136 576 -4080 610
rect -3820 576 -3764 610
rect -3504 576 -3448 610
rect -3188 576 -3132 610
rect -2872 576 -2816 610
rect -2556 576 -2500 610
rect -2240 576 -2184 610
rect -1924 576 -1868 610
rect -1608 576 -1552 610
rect -1292 576 -1236 610
rect -976 576 -920 610
rect -660 576 -604 610
rect -344 576 -288 610
rect -28 576 28 610
rect 288 576 344 610
rect 604 576 660 610
rect 920 576 976 610
rect 1236 576 1292 610
rect 1552 576 1608 610
rect 1868 576 1924 610
rect 2184 576 2240 610
rect 2500 576 2556 610
rect 2816 576 2872 610
rect 3132 576 3188 610
rect 3448 576 3504 610
rect 3764 576 3820 610
rect 4080 576 4136 610
rect 4396 576 4452 610
rect 4712 576 4768 610
rect 5028 576 5084 610
rect 5344 576 5400 610
rect 5660 576 5716 610
rect 5976 576 6032 610
rect 6292 576 6348 610
rect 6608 576 6664 610
rect 6924 576 6980 610
rect 7240 576 7296 610
rect 7556 576 7612 610
rect 7872 576 7928 610
rect 8188 576 8244 610
rect 8504 576 8560 610
rect 8820 576 8876 610
rect 9136 576 9192 610
rect 9452 576 9508 610
rect 9768 576 9824 610
rect 10084 576 10140 610
rect 10400 576 10456 610
rect 10716 576 10772 610
rect 11032 576 11088 610
rect 11348 576 11404 610
rect 11664 576 11720 610
rect 11980 576 12036 610
rect 12296 576 12352 610
rect 12612 576 12668 610
rect 12928 576 12984 610
rect -12984 567 -12928 576
rect -12668 567 -12612 576
rect -12352 567 -12296 576
rect -12036 567 -11980 576
rect -11720 567 -11664 576
rect -11404 567 -11348 576
rect -11088 567 -11032 576
rect -10772 567 -10716 576
rect -10456 567 -10400 576
rect -10140 567 -10084 576
rect -9824 567 -9768 576
rect -9508 567 -9452 576
rect -9192 567 -9136 576
rect -8876 567 -8820 576
rect -8560 567 -8504 576
rect -8244 567 -8188 576
rect -7928 567 -7872 576
rect -7612 567 -7556 576
rect -7296 567 -7240 576
rect -6980 567 -6924 576
rect -6664 567 -6608 576
rect -6348 567 -6292 576
rect -6032 567 -5976 576
rect -5716 567 -5660 576
rect -5400 567 -5344 576
rect -5084 567 -5028 576
rect -4768 567 -4712 576
rect -4452 567 -4396 576
rect -4136 567 -4080 576
rect -3820 567 -3764 576
rect -3504 567 -3448 576
rect -3188 567 -3132 576
rect -2872 567 -2816 576
rect -2556 567 -2500 576
rect -2240 567 -2184 576
rect -1924 567 -1868 576
rect -1608 567 -1552 576
rect -1292 567 -1236 576
rect -976 567 -920 576
rect -660 567 -604 576
rect -344 567 -288 576
rect -28 567 28 576
rect 288 567 344 576
rect 604 567 660 576
rect 920 567 976 576
rect 1236 567 1292 576
rect 1552 567 1608 576
rect 1868 567 1924 576
rect 2184 567 2240 576
rect 2500 567 2556 576
rect 2816 567 2872 576
rect 3132 567 3188 576
rect 3448 567 3504 576
rect 3764 567 3820 576
rect 4080 567 4136 576
rect 4396 567 4452 576
rect 4712 567 4768 576
rect 5028 567 5084 576
rect 5344 567 5400 576
rect 5660 567 5716 576
rect 5976 567 6032 576
rect 6292 567 6348 576
rect 6608 567 6664 576
rect 6924 567 6980 576
rect 7240 567 7296 576
rect 7556 567 7612 576
rect 7872 567 7928 576
rect 8188 567 8244 576
rect 8504 567 8560 576
rect 8820 567 8876 576
rect 9136 567 9192 576
rect 9452 567 9508 576
rect 9768 567 9824 576
rect 10084 567 10140 576
rect 10400 567 10456 576
rect 10716 567 10772 576
rect 11032 567 11088 576
rect 11348 567 11404 576
rect 11664 567 11720 576
rect 11980 567 12036 576
rect 12296 567 12352 576
rect 12612 567 12668 576
rect 12928 567 12984 576
rect -12982 388 -12930 394
rect -12982 -388 -12973 388
rect -12973 -388 -12939 388
rect -12939 -388 -12930 388
rect -12982 -394 -12930 -388
rect -12824 388 -12772 394
rect -12824 -388 -12815 388
rect -12815 -388 -12781 388
rect -12781 -388 -12772 388
rect -12824 -394 -12772 -388
rect -12666 388 -12614 394
rect -12666 -388 -12657 388
rect -12657 -388 -12623 388
rect -12623 -388 -12614 388
rect -12666 -394 -12614 -388
rect -12508 388 -12456 394
rect -12508 -388 -12499 388
rect -12499 -388 -12465 388
rect -12465 -388 -12456 388
rect -12508 -394 -12456 -388
rect -12350 388 -12298 394
rect -12350 -388 -12341 388
rect -12341 -388 -12307 388
rect -12307 -388 -12298 388
rect -12350 -394 -12298 -388
rect -12192 388 -12140 394
rect -12192 -388 -12183 388
rect -12183 -388 -12149 388
rect -12149 -388 -12140 388
rect -12192 -394 -12140 -388
rect -12034 388 -11982 394
rect -12034 -388 -12025 388
rect -12025 -388 -11991 388
rect -11991 -388 -11982 388
rect -12034 -394 -11982 -388
rect -11876 388 -11824 394
rect -11876 -388 -11867 388
rect -11867 -388 -11833 388
rect -11833 -388 -11824 388
rect -11876 -394 -11824 -388
rect -11718 388 -11666 394
rect -11718 -388 -11709 388
rect -11709 -388 -11675 388
rect -11675 -388 -11666 388
rect -11718 -394 -11666 -388
rect -11560 388 -11508 394
rect -11560 -388 -11551 388
rect -11551 -388 -11517 388
rect -11517 -388 -11508 388
rect -11560 -394 -11508 -388
rect -11402 388 -11350 394
rect -11402 -388 -11393 388
rect -11393 -388 -11359 388
rect -11359 -388 -11350 388
rect -11402 -394 -11350 -388
rect -11244 388 -11192 394
rect -11244 -388 -11235 388
rect -11235 -388 -11201 388
rect -11201 -388 -11192 388
rect -11244 -394 -11192 -388
rect -11086 388 -11034 394
rect -11086 -388 -11077 388
rect -11077 -388 -11043 388
rect -11043 -388 -11034 388
rect -11086 -394 -11034 -388
rect -10928 388 -10876 394
rect -10928 -388 -10919 388
rect -10919 -388 -10885 388
rect -10885 -388 -10876 388
rect -10928 -394 -10876 -388
rect -10770 388 -10718 394
rect -10770 -388 -10761 388
rect -10761 -388 -10727 388
rect -10727 -388 -10718 388
rect -10770 -394 -10718 -388
rect -10612 388 -10560 394
rect -10612 -388 -10603 388
rect -10603 -388 -10569 388
rect -10569 -388 -10560 388
rect -10612 -394 -10560 -388
rect -10454 388 -10402 394
rect -10454 -388 -10445 388
rect -10445 -388 -10411 388
rect -10411 -388 -10402 388
rect -10454 -394 -10402 -388
rect -10296 388 -10244 394
rect -10296 -388 -10287 388
rect -10287 -388 -10253 388
rect -10253 -388 -10244 388
rect -10296 -394 -10244 -388
rect -10138 388 -10086 394
rect -10138 -388 -10129 388
rect -10129 -388 -10095 388
rect -10095 -388 -10086 388
rect -10138 -394 -10086 -388
rect -9980 388 -9928 394
rect -9980 -388 -9971 388
rect -9971 -388 -9937 388
rect -9937 -388 -9928 388
rect -9980 -394 -9928 -388
rect -9822 388 -9770 394
rect -9822 -388 -9813 388
rect -9813 -388 -9779 388
rect -9779 -388 -9770 388
rect -9822 -394 -9770 -388
rect -9664 388 -9612 394
rect -9664 -388 -9655 388
rect -9655 -388 -9621 388
rect -9621 -388 -9612 388
rect -9664 -394 -9612 -388
rect -9506 388 -9454 394
rect -9506 -388 -9497 388
rect -9497 -388 -9463 388
rect -9463 -388 -9454 388
rect -9506 -394 -9454 -388
rect -9348 388 -9296 394
rect -9348 -388 -9339 388
rect -9339 -388 -9305 388
rect -9305 -388 -9296 388
rect -9348 -394 -9296 -388
rect -9190 388 -9138 394
rect -9190 -388 -9181 388
rect -9181 -388 -9147 388
rect -9147 -388 -9138 388
rect -9190 -394 -9138 -388
rect -9032 388 -8980 394
rect -9032 -388 -9023 388
rect -9023 -388 -8989 388
rect -8989 -388 -8980 388
rect -9032 -394 -8980 -388
rect -8874 388 -8822 394
rect -8874 -388 -8865 388
rect -8865 -388 -8831 388
rect -8831 -388 -8822 388
rect -8874 -394 -8822 -388
rect -8716 388 -8664 394
rect -8716 -388 -8707 388
rect -8707 -388 -8673 388
rect -8673 -388 -8664 388
rect -8716 -394 -8664 -388
rect -8558 388 -8506 394
rect -8558 -388 -8549 388
rect -8549 -388 -8515 388
rect -8515 -388 -8506 388
rect -8558 -394 -8506 -388
rect -8400 388 -8348 394
rect -8400 -388 -8391 388
rect -8391 -388 -8357 388
rect -8357 -388 -8348 388
rect -8400 -394 -8348 -388
rect -8242 388 -8190 394
rect -8242 -388 -8233 388
rect -8233 -388 -8199 388
rect -8199 -388 -8190 388
rect -8242 -394 -8190 -388
rect -8084 388 -8032 394
rect -8084 -388 -8075 388
rect -8075 -388 -8041 388
rect -8041 -388 -8032 388
rect -8084 -394 -8032 -388
rect -7926 388 -7874 394
rect -7926 -388 -7917 388
rect -7917 -388 -7883 388
rect -7883 -388 -7874 388
rect -7926 -394 -7874 -388
rect -7768 388 -7716 394
rect -7768 -388 -7759 388
rect -7759 -388 -7725 388
rect -7725 -388 -7716 388
rect -7768 -394 -7716 -388
rect -7610 388 -7558 394
rect -7610 -388 -7601 388
rect -7601 -388 -7567 388
rect -7567 -388 -7558 388
rect -7610 -394 -7558 -388
rect -7452 388 -7400 394
rect -7452 -388 -7443 388
rect -7443 -388 -7409 388
rect -7409 -388 -7400 388
rect -7452 -394 -7400 -388
rect -7294 388 -7242 394
rect -7294 -388 -7285 388
rect -7285 -388 -7251 388
rect -7251 -388 -7242 388
rect -7294 -394 -7242 -388
rect -7136 388 -7084 394
rect -7136 -388 -7127 388
rect -7127 -388 -7093 388
rect -7093 -388 -7084 388
rect -7136 -394 -7084 -388
rect -6978 388 -6926 394
rect -6978 -388 -6969 388
rect -6969 -388 -6935 388
rect -6935 -388 -6926 388
rect -6978 -394 -6926 -388
rect -6820 388 -6768 394
rect -6820 -388 -6811 388
rect -6811 -388 -6777 388
rect -6777 -388 -6768 388
rect -6820 -394 -6768 -388
rect -6662 388 -6610 394
rect -6662 -388 -6653 388
rect -6653 -388 -6619 388
rect -6619 -388 -6610 388
rect -6662 -394 -6610 -388
rect -6504 388 -6452 394
rect -6504 -388 -6495 388
rect -6495 -388 -6461 388
rect -6461 -388 -6452 388
rect -6504 -394 -6452 -388
rect -6346 388 -6294 394
rect -6346 -388 -6337 388
rect -6337 -388 -6303 388
rect -6303 -388 -6294 388
rect -6346 -394 -6294 -388
rect -6188 388 -6136 394
rect -6188 -388 -6179 388
rect -6179 -388 -6145 388
rect -6145 -388 -6136 388
rect -6188 -394 -6136 -388
rect -6030 388 -5978 394
rect -6030 -388 -6021 388
rect -6021 -388 -5987 388
rect -5987 -388 -5978 388
rect -6030 -394 -5978 -388
rect -5872 388 -5820 394
rect -5872 -388 -5863 388
rect -5863 -388 -5829 388
rect -5829 -388 -5820 388
rect -5872 -394 -5820 -388
rect -5714 388 -5662 394
rect -5714 -388 -5705 388
rect -5705 -388 -5671 388
rect -5671 -388 -5662 388
rect -5714 -394 -5662 -388
rect -5556 388 -5504 394
rect -5556 -388 -5547 388
rect -5547 -388 -5513 388
rect -5513 -388 -5504 388
rect -5556 -394 -5504 -388
rect -5398 388 -5346 394
rect -5398 -388 -5389 388
rect -5389 -388 -5355 388
rect -5355 -388 -5346 388
rect -5398 -394 -5346 -388
rect -5240 388 -5188 394
rect -5240 -388 -5231 388
rect -5231 -388 -5197 388
rect -5197 -388 -5188 388
rect -5240 -394 -5188 -388
rect -5082 388 -5030 394
rect -5082 -388 -5073 388
rect -5073 -388 -5039 388
rect -5039 -388 -5030 388
rect -5082 -394 -5030 -388
rect -4924 388 -4872 394
rect -4924 -388 -4915 388
rect -4915 -388 -4881 388
rect -4881 -388 -4872 388
rect -4924 -394 -4872 -388
rect -4766 388 -4714 394
rect -4766 -388 -4757 388
rect -4757 -388 -4723 388
rect -4723 -388 -4714 388
rect -4766 -394 -4714 -388
rect -4450 388 -4398 394
rect -4450 -388 -4441 388
rect -4441 -388 -4407 388
rect -4407 -388 -4398 388
rect -4450 -394 -4398 -388
rect -4292 388 -4240 394
rect -4292 -388 -4283 388
rect -4283 -388 -4249 388
rect -4249 -388 -4240 388
rect -4292 -394 -4240 -388
rect -4134 388 -4082 394
rect -4134 -388 -4125 388
rect -4125 -388 -4091 388
rect -4091 -388 -4082 388
rect -4134 -394 -4082 -388
rect -3976 388 -3924 394
rect -3976 -388 -3967 388
rect -3967 -388 -3933 388
rect -3933 -388 -3924 388
rect -3976 -394 -3924 -388
rect -3818 388 -3766 394
rect -3818 -388 -3809 388
rect -3809 -388 -3775 388
rect -3775 -388 -3766 388
rect -3818 -394 -3766 -388
rect -3660 388 -3608 394
rect -3660 -388 -3651 388
rect -3651 -388 -3617 388
rect -3617 -388 -3608 388
rect -3660 -394 -3608 -388
rect -3502 388 -3450 394
rect -3502 -388 -3493 388
rect -3493 -388 -3459 388
rect -3459 -388 -3450 388
rect -3502 -394 -3450 -388
rect -3344 388 -3292 394
rect -3344 -388 -3335 388
rect -3335 -388 -3301 388
rect -3301 -388 -3292 388
rect -3344 -394 -3292 -388
rect -3186 388 -3134 394
rect -3186 -388 -3177 388
rect -3177 -388 -3143 388
rect -3143 -388 -3134 388
rect -3186 -394 -3134 -388
rect -3028 388 -2976 394
rect -3028 -388 -3019 388
rect -3019 -388 -2985 388
rect -2985 -388 -2976 388
rect -3028 -394 -2976 -388
rect -2870 388 -2818 394
rect -2870 -388 -2861 388
rect -2861 -388 -2827 388
rect -2827 -388 -2818 388
rect -2870 -394 -2818 -388
rect -2712 388 -2660 394
rect -2712 -388 -2703 388
rect -2703 -388 -2669 388
rect -2669 -388 -2660 388
rect -2712 -394 -2660 -388
rect -2554 388 -2502 394
rect -2554 -388 -2545 388
rect -2545 -388 -2511 388
rect -2511 -388 -2502 388
rect -2554 -394 -2502 -388
rect -2396 388 -2344 394
rect -2396 -388 -2387 388
rect -2387 -388 -2353 388
rect -2353 -388 -2344 388
rect -2396 -394 -2344 -388
rect -2238 388 -2186 394
rect -2238 -388 -2229 388
rect -2229 -388 -2195 388
rect -2195 -388 -2186 388
rect -2238 -394 -2186 -388
rect -2080 388 -2028 394
rect -2080 -388 -2071 388
rect -2071 -388 -2037 388
rect -2037 -388 -2028 388
rect -2080 -394 -2028 -388
rect -1922 388 -1870 394
rect -1922 -388 -1913 388
rect -1913 -388 -1879 388
rect -1879 -388 -1870 388
rect -1922 -394 -1870 -388
rect -1764 388 -1712 394
rect -1764 -388 -1755 388
rect -1755 -388 -1721 388
rect -1721 -388 -1712 388
rect -1764 -394 -1712 -388
rect -1606 388 -1554 394
rect -1606 -388 -1597 388
rect -1597 -388 -1563 388
rect -1563 -388 -1554 388
rect -1606 -394 -1554 -388
rect -1448 388 -1396 394
rect -1448 -388 -1439 388
rect -1439 -388 -1405 388
rect -1405 -388 -1396 388
rect -1448 -394 -1396 -388
rect -1290 388 -1238 394
rect -1290 -388 -1281 388
rect -1281 -388 -1247 388
rect -1247 -388 -1238 388
rect -1290 -394 -1238 -388
rect -1132 388 -1080 394
rect -1132 -388 -1123 388
rect -1123 -388 -1089 388
rect -1089 -388 -1080 388
rect -1132 -394 -1080 -388
rect -974 388 -922 394
rect -974 -388 -965 388
rect -965 -388 -931 388
rect -931 -388 -922 388
rect -974 -394 -922 -388
rect -816 388 -764 394
rect -816 -388 -807 388
rect -807 -388 -773 388
rect -773 -388 -764 388
rect -816 -394 -764 -388
rect -658 388 -606 394
rect -658 -388 -649 388
rect -649 -388 -615 388
rect -615 -388 -606 388
rect -658 -394 -606 -388
rect -500 388 -448 394
rect -500 -388 -491 388
rect -491 -388 -457 388
rect -457 -388 -448 388
rect -500 -394 -448 -388
rect -342 388 -290 394
rect -342 -388 -333 388
rect -333 -388 -299 388
rect -299 -388 -290 388
rect -342 -394 -290 -388
rect -184 388 -132 394
rect -184 -388 -175 388
rect -175 -388 -141 388
rect -141 -388 -132 388
rect -184 -394 -132 -388
rect -26 388 26 394
rect -26 -388 -17 388
rect -17 -388 17 388
rect 17 -388 26 388
rect -26 -394 26 -388
rect 132 388 184 394
rect 132 -388 141 388
rect 141 -388 175 388
rect 175 -388 184 388
rect 132 -394 184 -388
rect 290 388 342 394
rect 290 -388 299 388
rect 299 -388 333 388
rect 333 -388 342 388
rect 290 -394 342 -388
rect 448 388 500 394
rect 448 -388 457 388
rect 457 -388 491 388
rect 491 -388 500 388
rect 448 -394 500 -388
rect 606 388 658 394
rect 606 -388 615 388
rect 615 -388 649 388
rect 649 -388 658 388
rect 606 -394 658 -388
rect 764 388 816 394
rect 764 -388 773 388
rect 773 -388 807 388
rect 807 -388 816 388
rect 764 -394 816 -388
rect 922 388 974 394
rect 922 -388 931 388
rect 931 -388 965 388
rect 965 -388 974 388
rect 922 -394 974 -388
rect 1080 388 1132 394
rect 1080 -388 1089 388
rect 1089 -388 1123 388
rect 1123 -388 1132 388
rect 1080 -394 1132 -388
rect 1238 388 1290 394
rect 1238 -388 1247 388
rect 1247 -388 1281 388
rect 1281 -388 1290 388
rect 1238 -394 1290 -388
rect 1396 388 1448 394
rect 1396 -388 1405 388
rect 1405 -388 1439 388
rect 1439 -388 1448 388
rect 1396 -394 1448 -388
rect 1554 388 1606 394
rect 1554 -388 1563 388
rect 1563 -388 1597 388
rect 1597 -388 1606 388
rect 1554 -394 1606 -388
rect 1712 388 1764 394
rect 1712 -388 1721 388
rect 1721 -388 1755 388
rect 1755 -388 1764 388
rect 1712 -394 1764 -388
rect 1870 388 1922 394
rect 1870 -388 1879 388
rect 1879 -388 1913 388
rect 1913 -388 1922 388
rect 1870 -394 1922 -388
rect 2028 388 2080 394
rect 2028 -388 2037 388
rect 2037 -388 2071 388
rect 2071 -388 2080 388
rect 2028 -394 2080 -388
rect 2186 388 2238 394
rect 2186 -388 2195 388
rect 2195 -388 2229 388
rect 2229 -388 2238 388
rect 2186 -394 2238 -388
rect 2344 388 2396 394
rect 2344 -388 2353 388
rect 2353 -388 2387 388
rect 2387 -388 2396 388
rect 2344 -394 2396 -388
rect 2502 388 2554 394
rect 2502 -388 2511 388
rect 2511 -388 2545 388
rect 2545 -388 2554 388
rect 2502 -394 2554 -388
rect 2660 388 2712 394
rect 2660 -388 2669 388
rect 2669 -388 2703 388
rect 2703 -388 2712 388
rect 2660 -394 2712 -388
rect 2818 388 2870 394
rect 2818 -388 2827 388
rect 2827 -388 2861 388
rect 2861 -388 2870 388
rect 2818 -394 2870 -388
rect 2976 388 3028 394
rect 2976 -388 2985 388
rect 2985 -388 3019 388
rect 3019 -388 3028 388
rect 2976 -394 3028 -388
rect 3134 388 3186 394
rect 3134 -388 3143 388
rect 3143 -388 3177 388
rect 3177 -388 3186 388
rect 3134 -394 3186 -388
rect 3292 388 3344 394
rect 3292 -388 3301 388
rect 3301 -388 3335 388
rect 3335 -388 3344 388
rect 3292 -394 3344 -388
rect 3450 388 3502 394
rect 3450 -388 3459 388
rect 3459 -388 3493 388
rect 3493 -388 3502 388
rect 3450 -394 3502 -388
rect 3608 388 3660 394
rect 3608 -388 3617 388
rect 3617 -388 3651 388
rect 3651 -388 3660 388
rect 3608 -394 3660 -388
rect 3766 388 3818 394
rect 3766 -388 3775 388
rect 3775 -388 3809 388
rect 3809 -388 3818 388
rect 3766 -394 3818 -388
rect 3924 388 3976 394
rect 3924 -388 3933 388
rect 3933 -388 3967 388
rect 3967 -388 3976 388
rect 3924 -394 3976 -388
rect 4082 388 4134 394
rect 4082 -388 4091 388
rect 4091 -388 4125 388
rect 4125 -388 4134 388
rect 4082 -394 4134 -388
rect 4240 388 4292 394
rect 4240 -388 4249 388
rect 4249 -388 4283 388
rect 4283 -388 4292 388
rect 4240 -394 4292 -388
rect 4398 388 4450 394
rect 4398 -388 4407 388
rect 4407 -388 4441 388
rect 4441 -388 4450 388
rect 4398 -394 4450 -388
rect 4714 388 4766 394
rect 4714 -388 4723 388
rect 4723 -388 4757 388
rect 4757 -388 4766 388
rect 4714 -394 4766 -388
rect 4872 388 4924 394
rect 4872 -388 4881 388
rect 4881 -388 4915 388
rect 4915 -388 4924 388
rect 4872 -394 4924 -388
rect 5030 388 5082 394
rect 5030 -388 5039 388
rect 5039 -388 5073 388
rect 5073 -388 5082 388
rect 5030 -394 5082 -388
rect 5188 388 5240 394
rect 5188 -388 5197 388
rect 5197 -388 5231 388
rect 5231 -388 5240 388
rect 5188 -394 5240 -388
rect 5346 388 5398 394
rect 5346 -388 5355 388
rect 5355 -388 5389 388
rect 5389 -388 5398 388
rect 5346 -394 5398 -388
rect 5504 388 5556 394
rect 5504 -388 5513 388
rect 5513 -388 5547 388
rect 5547 -388 5556 388
rect 5504 -394 5556 -388
rect 5662 388 5714 394
rect 5662 -388 5671 388
rect 5671 -388 5705 388
rect 5705 -388 5714 388
rect 5662 -394 5714 -388
rect 5820 388 5872 394
rect 5820 -388 5829 388
rect 5829 -388 5863 388
rect 5863 -388 5872 388
rect 5820 -394 5872 -388
rect 5978 388 6030 394
rect 5978 -388 5987 388
rect 5987 -388 6021 388
rect 6021 -388 6030 388
rect 5978 -394 6030 -388
rect 6136 388 6188 394
rect 6136 -388 6145 388
rect 6145 -388 6179 388
rect 6179 -388 6188 388
rect 6136 -394 6188 -388
rect 6294 388 6346 394
rect 6294 -388 6303 388
rect 6303 -388 6337 388
rect 6337 -388 6346 388
rect 6294 -394 6346 -388
rect 6452 388 6504 394
rect 6452 -388 6461 388
rect 6461 -388 6495 388
rect 6495 -388 6504 388
rect 6452 -394 6504 -388
rect 6610 388 6662 394
rect 6610 -388 6619 388
rect 6619 -388 6653 388
rect 6653 -388 6662 388
rect 6610 -394 6662 -388
rect 6768 388 6820 394
rect 6768 -388 6777 388
rect 6777 -388 6811 388
rect 6811 -388 6820 388
rect 6768 -394 6820 -388
rect 6926 388 6978 394
rect 6926 -388 6935 388
rect 6935 -388 6969 388
rect 6969 -388 6978 388
rect 6926 -394 6978 -388
rect 7084 388 7136 394
rect 7084 -388 7093 388
rect 7093 -388 7127 388
rect 7127 -388 7136 388
rect 7084 -394 7136 -388
rect 7242 388 7294 394
rect 7242 -388 7251 388
rect 7251 -388 7285 388
rect 7285 -388 7294 388
rect 7242 -394 7294 -388
rect 7400 388 7452 394
rect 7400 -388 7409 388
rect 7409 -388 7443 388
rect 7443 -388 7452 388
rect 7400 -394 7452 -388
rect 7558 388 7610 394
rect 7558 -388 7567 388
rect 7567 -388 7601 388
rect 7601 -388 7610 388
rect 7558 -394 7610 -388
rect 7716 388 7768 394
rect 7716 -388 7725 388
rect 7725 -388 7759 388
rect 7759 -388 7768 388
rect 7716 -394 7768 -388
rect 7874 388 7926 394
rect 7874 -388 7883 388
rect 7883 -388 7917 388
rect 7917 -388 7926 388
rect 7874 -394 7926 -388
rect 8032 388 8084 394
rect 8032 -388 8041 388
rect 8041 -388 8075 388
rect 8075 -388 8084 388
rect 8032 -394 8084 -388
rect 8190 388 8242 394
rect 8190 -388 8199 388
rect 8199 -388 8233 388
rect 8233 -388 8242 388
rect 8190 -394 8242 -388
rect 8348 388 8400 394
rect 8348 -388 8357 388
rect 8357 -388 8391 388
rect 8391 -388 8400 388
rect 8348 -394 8400 -388
rect 8506 388 8558 394
rect 8506 -388 8515 388
rect 8515 -388 8549 388
rect 8549 -388 8558 388
rect 8506 -394 8558 -388
rect 8664 388 8716 394
rect 8664 -388 8673 388
rect 8673 -388 8707 388
rect 8707 -388 8716 388
rect 8664 -394 8716 -388
rect 8822 388 8874 394
rect 8822 -388 8831 388
rect 8831 -388 8865 388
rect 8865 -388 8874 388
rect 8822 -394 8874 -388
rect 8980 388 9032 394
rect 8980 -388 8989 388
rect 8989 -388 9023 388
rect 9023 -388 9032 388
rect 8980 -394 9032 -388
rect 9138 388 9190 394
rect 9138 -388 9147 388
rect 9147 -388 9181 388
rect 9181 -388 9190 388
rect 9138 -394 9190 -388
rect 9296 388 9348 394
rect 9296 -388 9305 388
rect 9305 -388 9339 388
rect 9339 -388 9348 388
rect 9296 -394 9348 -388
rect 9454 388 9506 394
rect 9454 -388 9463 388
rect 9463 -388 9497 388
rect 9497 -388 9506 388
rect 9454 -394 9506 -388
rect 9612 388 9664 394
rect 9612 -388 9621 388
rect 9621 -388 9655 388
rect 9655 -388 9664 388
rect 9612 -394 9664 -388
rect 9770 388 9822 394
rect 9770 -388 9779 388
rect 9779 -388 9813 388
rect 9813 -388 9822 388
rect 9770 -394 9822 -388
rect 9928 388 9980 394
rect 9928 -388 9937 388
rect 9937 -388 9971 388
rect 9971 -388 9980 388
rect 9928 -394 9980 -388
rect 10086 388 10138 394
rect 10086 -388 10095 388
rect 10095 -388 10129 388
rect 10129 -388 10138 388
rect 10086 -394 10138 -388
rect 10244 388 10296 394
rect 10244 -388 10253 388
rect 10253 -388 10287 388
rect 10287 -388 10296 388
rect 10244 -394 10296 -388
rect 10402 388 10454 394
rect 10402 -388 10411 388
rect 10411 -388 10445 388
rect 10445 -388 10454 388
rect 10402 -394 10454 -388
rect 10560 388 10612 394
rect 10560 -388 10569 388
rect 10569 -388 10603 388
rect 10603 -388 10612 388
rect 10560 -394 10612 -388
rect 10718 388 10770 394
rect 10718 -388 10727 388
rect 10727 -388 10761 388
rect 10761 -388 10770 388
rect 10718 -394 10770 -388
rect 10876 388 10928 394
rect 10876 -388 10885 388
rect 10885 -388 10919 388
rect 10919 -388 10928 388
rect 10876 -394 10928 -388
rect 11034 388 11086 394
rect 11034 -388 11043 388
rect 11043 -388 11077 388
rect 11077 -388 11086 388
rect 11034 -394 11086 -388
rect 11192 388 11244 394
rect 11192 -388 11201 388
rect 11201 -388 11235 388
rect 11235 -388 11244 388
rect 11192 -394 11244 -388
rect 11350 388 11402 394
rect 11350 -388 11359 388
rect 11359 -388 11393 388
rect 11393 -388 11402 388
rect 11350 -394 11402 -388
rect 11508 388 11560 394
rect 11508 -388 11517 388
rect 11517 -388 11551 388
rect 11551 -388 11560 388
rect 11508 -394 11560 -388
rect 11666 388 11718 394
rect 11666 -388 11675 388
rect 11675 -388 11709 388
rect 11709 -388 11718 388
rect 11666 -394 11718 -388
rect 11824 388 11876 394
rect 11824 -388 11833 388
rect 11833 -388 11867 388
rect 11867 -388 11876 388
rect 11824 -394 11876 -388
rect 11982 388 12034 394
rect 11982 -388 11991 388
rect 11991 -388 12025 388
rect 12025 -388 12034 388
rect 11982 -394 12034 -388
rect 12140 388 12192 394
rect 12140 -388 12149 388
rect 12149 -388 12183 388
rect 12183 -388 12192 388
rect 12140 -394 12192 -388
rect 12298 388 12350 394
rect 12298 -388 12307 388
rect 12307 -388 12341 388
rect 12341 -388 12350 388
rect 12298 -394 12350 -388
rect 12456 388 12508 394
rect 12456 -388 12465 388
rect 12465 -388 12499 388
rect 12499 -388 12508 388
rect 12456 -394 12508 -388
rect 12614 388 12666 394
rect 12614 -388 12623 388
rect 12623 -388 12657 388
rect 12657 -388 12666 388
rect 12614 -394 12666 -388
rect 12772 388 12824 394
rect 12772 -388 12781 388
rect 12781 -388 12815 388
rect 12815 -388 12824 388
rect 12772 -394 12824 -388
rect 12930 388 12982 394
rect 12930 -388 12939 388
rect 12939 -388 12973 388
rect 12973 -388 12982 388
rect 12930 -394 12982 -388
rect -12984 -576 -12928 -567
rect -12668 -576 -12612 -567
rect -12352 -576 -12296 -567
rect -12036 -576 -11980 -567
rect -11720 -576 -11664 -567
rect -11404 -576 -11348 -567
rect -11088 -576 -11032 -567
rect -10772 -576 -10716 -567
rect -10456 -576 -10400 -567
rect -10140 -576 -10084 -567
rect -9824 -576 -9768 -567
rect -9508 -576 -9452 -567
rect -9192 -576 -9136 -567
rect -8876 -576 -8820 -567
rect -8560 -576 -8504 -567
rect -8244 -576 -8188 -567
rect -7928 -576 -7872 -567
rect -7612 -576 -7556 -567
rect -7296 -576 -7240 -567
rect -6980 -576 -6924 -567
rect -6664 -576 -6608 -567
rect -6348 -576 -6292 -567
rect -6032 -576 -5976 -567
rect -5716 -576 -5660 -567
rect -5400 -576 -5344 -567
rect -5084 -576 -5028 -567
rect -4768 -576 -4712 -567
rect -4452 -576 -4396 -567
rect -4136 -576 -4080 -567
rect -3820 -576 -3764 -567
rect -3504 -576 -3448 -567
rect -3188 -576 -3132 -567
rect -2872 -576 -2816 -567
rect -2556 -576 -2500 -567
rect -2240 -576 -2184 -567
rect -1924 -576 -1868 -567
rect -1608 -576 -1552 -567
rect -1292 -576 -1236 -567
rect -976 -576 -920 -567
rect -660 -576 -604 -567
rect -344 -576 -288 -567
rect -28 -576 28 -567
rect 288 -576 344 -567
rect 604 -576 660 -567
rect 920 -576 976 -567
rect 1236 -576 1292 -567
rect 1552 -576 1608 -567
rect 1868 -576 1924 -567
rect 2184 -576 2240 -567
rect 2500 -576 2556 -567
rect 2816 -576 2872 -567
rect 3132 -576 3188 -567
rect 3448 -576 3504 -567
rect 3764 -576 3820 -567
rect 4080 -576 4136 -567
rect 4396 -576 4452 -567
rect 4712 -576 4768 -567
rect 5028 -576 5084 -567
rect 5344 -576 5400 -567
rect 5660 -576 5716 -567
rect 5976 -576 6032 -567
rect 6292 -576 6348 -567
rect 6608 -576 6664 -567
rect 6924 -576 6980 -567
rect 7240 -576 7296 -567
rect 7556 -576 7612 -567
rect 7872 -576 7928 -567
rect 8188 -576 8244 -567
rect 8504 -576 8560 -567
rect 8820 -576 8876 -567
rect 9136 -576 9192 -567
rect 9452 -576 9508 -567
rect 9768 -576 9824 -567
rect 10084 -576 10140 -567
rect 10400 -576 10456 -567
rect 10716 -576 10772 -567
rect 11032 -576 11088 -567
rect 11348 -576 11404 -567
rect 11664 -576 11720 -567
rect 11980 -576 12036 -567
rect 12296 -576 12352 -567
rect 12612 -576 12668 -567
rect 12928 -576 12984 -567
rect -12984 -610 -12928 -576
rect -12668 -610 -12612 -576
rect -12352 -610 -12296 -576
rect -12036 -610 -11980 -576
rect -11720 -610 -11664 -576
rect -11404 -610 -11348 -576
rect -11088 -610 -11032 -576
rect -10772 -610 -10716 -576
rect -10456 -610 -10400 -576
rect -10140 -610 -10084 -576
rect -9824 -610 -9768 -576
rect -9508 -610 -9452 -576
rect -9192 -610 -9136 -576
rect -8876 -610 -8820 -576
rect -8560 -610 -8504 -576
rect -8244 -610 -8188 -576
rect -7928 -610 -7872 -576
rect -7612 -610 -7556 -576
rect -7296 -610 -7240 -576
rect -6980 -610 -6924 -576
rect -6664 -610 -6608 -576
rect -6348 -610 -6292 -576
rect -6032 -610 -5976 -576
rect -5716 -610 -5660 -576
rect -5400 -610 -5344 -576
rect -5084 -610 -5028 -576
rect -4768 -610 -4712 -576
rect -4452 -610 -4396 -576
rect -4136 -610 -4080 -576
rect -3820 -610 -3764 -576
rect -3504 -610 -3448 -576
rect -3188 -610 -3132 -576
rect -2872 -610 -2816 -576
rect -2556 -610 -2500 -576
rect -2240 -610 -2184 -576
rect -1924 -610 -1868 -576
rect -1608 -610 -1552 -576
rect -1292 -610 -1236 -576
rect -976 -610 -920 -576
rect -660 -610 -604 -576
rect -344 -610 -288 -576
rect -28 -610 28 -576
rect 288 -610 344 -576
rect 604 -610 660 -576
rect 920 -610 976 -576
rect 1236 -610 1292 -576
rect 1552 -610 1608 -576
rect 1868 -610 1924 -576
rect 2184 -610 2240 -576
rect 2500 -610 2556 -576
rect 2816 -610 2872 -576
rect 3132 -610 3188 -576
rect 3448 -610 3504 -576
rect 3764 -610 3820 -576
rect 4080 -610 4136 -576
rect 4396 -610 4452 -576
rect 4712 -610 4768 -576
rect 5028 -610 5084 -576
rect 5344 -610 5400 -576
rect 5660 -610 5716 -576
rect 5976 -610 6032 -576
rect 6292 -610 6348 -576
rect 6608 -610 6664 -576
rect 6924 -610 6980 -576
rect 7240 -610 7296 -576
rect 7556 -610 7612 -576
rect 7872 -610 7928 -576
rect 8188 -610 8244 -576
rect 8504 -610 8560 -576
rect 8820 -610 8876 -576
rect 9136 -610 9192 -576
rect 9452 -610 9508 -576
rect 9768 -610 9824 -576
rect 10084 -610 10140 -576
rect 10400 -610 10456 -576
rect 10716 -610 10772 -576
rect 11032 -610 11088 -576
rect 11348 -610 11404 -576
rect 11664 -610 11720 -576
rect 11980 -610 12036 -576
rect 12296 -610 12352 -576
rect 12612 -610 12668 -576
rect 12928 -610 12984 -576
rect -12984 -619 -12928 -610
rect -12668 -619 -12612 -610
rect -12352 -619 -12296 -610
rect -12036 -619 -11980 -610
rect -11720 -619 -11664 -610
rect -11404 -619 -11348 -610
rect -11088 -619 -11032 -610
rect -10772 -619 -10716 -610
rect -10456 -619 -10400 -610
rect -10140 -619 -10084 -610
rect -9824 -619 -9768 -610
rect -9508 -619 -9452 -610
rect -9192 -619 -9136 -610
rect -8876 -619 -8820 -610
rect -8560 -619 -8504 -610
rect -8244 -619 -8188 -610
rect -7928 -619 -7872 -610
rect -7612 -619 -7556 -610
rect -7296 -619 -7240 -610
rect -6980 -619 -6924 -610
rect -6664 -619 -6608 -610
rect -6348 -619 -6292 -610
rect -6032 -619 -5976 -610
rect -5716 -619 -5660 -610
rect -5400 -619 -5344 -610
rect -5084 -619 -5028 -610
rect -4768 -619 -4712 -610
rect -4452 -619 -4396 -610
rect -4136 -619 -4080 -610
rect -3820 -619 -3764 -610
rect -3504 -619 -3448 -610
rect -3188 -619 -3132 -610
rect -2872 -619 -2816 -610
rect -2556 -619 -2500 -610
rect -2240 -619 -2184 -610
rect -1924 -619 -1868 -610
rect -1608 -619 -1552 -610
rect -1292 -619 -1236 -610
rect -976 -619 -920 -610
rect -660 -619 -604 -610
rect -344 -619 -288 -610
rect -28 -619 28 -610
rect 288 -619 344 -610
rect 604 -619 660 -610
rect 920 -619 976 -610
rect 1236 -619 1292 -610
rect 1552 -619 1608 -610
rect 1868 -619 1924 -610
rect 2184 -619 2240 -610
rect 2500 -619 2556 -610
rect 2816 -619 2872 -610
rect 3132 -619 3188 -610
rect 3448 -619 3504 -610
rect 3764 -619 3820 -610
rect 4080 -619 4136 -610
rect 4396 -619 4452 -610
rect 4712 -619 4768 -610
rect 5028 -619 5084 -610
rect 5344 -619 5400 -610
rect 5660 -619 5716 -610
rect 5976 -619 6032 -610
rect 6292 -619 6348 -610
rect 6608 -619 6664 -610
rect 6924 -619 6980 -610
rect 7240 -619 7296 -610
rect 7556 -619 7612 -610
rect 7872 -619 7928 -610
rect 8188 -619 8244 -610
rect 8504 -619 8560 -610
rect 8820 -619 8876 -610
rect 9136 -619 9192 -610
rect 9452 -619 9508 -610
rect 9768 -619 9824 -610
rect 10084 -619 10140 -610
rect 10400 -619 10456 -610
rect 10716 -619 10772 -610
rect 11032 -619 11088 -610
rect 11348 -619 11404 -610
rect 11664 -619 11720 -610
rect 11980 -619 12036 -610
rect 12296 -619 12352 -610
rect 12612 -619 12668 -610
rect 12928 -619 12984 -610
<< metal2 >>
rect -12984 619 -12928 700
rect -12984 394 -12928 567
rect -12984 295 -12982 394
rect -12930 295 -12928 394
rect -12984 -394 -12982 -295
rect -12930 -394 -12928 -295
rect -12984 -567 -12928 -394
rect -12984 -700 -12928 -619
rect -12826 394 -12770 700
rect -12826 -385 -12824 394
rect -12772 -385 -12770 394
rect -12826 -700 -12770 -691
rect -12668 619 -12612 700
rect -12668 394 -12612 567
rect -12668 295 -12666 394
rect -12614 295 -12612 394
rect -12668 -394 -12666 -295
rect -12614 -394 -12612 -295
rect -12668 -567 -12612 -394
rect -12668 -700 -12612 -619
rect -12510 691 -12454 700
rect -12510 -394 -12508 385
rect -12456 -394 -12454 385
rect -12510 -700 -12454 -394
rect -12352 619 -12296 700
rect -12352 394 -12296 567
rect -12352 295 -12350 394
rect -12298 295 -12296 394
rect -12352 -394 -12350 -295
rect -12298 -394 -12296 -295
rect -12352 -567 -12296 -394
rect -12352 -700 -12296 -619
rect -12194 394 -12138 700
rect -12194 -385 -12192 394
rect -12140 -385 -12138 394
rect -12194 -700 -12138 -691
rect -12036 619 -11980 700
rect -12036 394 -11980 567
rect -12036 295 -12034 394
rect -11982 295 -11980 394
rect -12036 -394 -12034 -295
rect -11982 -394 -11980 -295
rect -12036 -567 -11980 -394
rect -12036 -700 -11980 -619
rect -11878 691 -11822 700
rect -11878 -394 -11876 385
rect -11824 -394 -11822 385
rect -11878 -700 -11822 -394
rect -11720 619 -11664 700
rect -11720 394 -11664 567
rect -11720 295 -11718 394
rect -11666 295 -11664 394
rect -11720 -394 -11718 -295
rect -11666 -394 -11664 -295
rect -11720 -567 -11664 -394
rect -11720 -700 -11664 -619
rect -11562 394 -11506 700
rect -11562 -385 -11560 394
rect -11508 -385 -11506 394
rect -11562 -700 -11506 -691
rect -11404 619 -11348 700
rect -11404 394 -11348 567
rect -11404 295 -11402 394
rect -11350 295 -11348 394
rect -11404 -394 -11402 -295
rect -11350 -394 -11348 -295
rect -11404 -567 -11348 -394
rect -11404 -700 -11348 -619
rect -11246 691 -11190 700
rect -11246 -394 -11244 385
rect -11192 -394 -11190 385
rect -11246 -700 -11190 -394
rect -11088 619 -11032 700
rect -11088 394 -11032 567
rect -11088 295 -11086 394
rect -11034 295 -11032 394
rect -11088 -394 -11086 -295
rect -11034 -394 -11032 -295
rect -11088 -567 -11032 -394
rect -11088 -700 -11032 -619
rect -10930 394 -10874 700
rect -10930 -385 -10928 394
rect -10876 -385 -10874 394
rect -10930 -700 -10874 -691
rect -10772 619 -10716 700
rect -10772 394 -10716 567
rect -10772 295 -10770 394
rect -10718 295 -10716 394
rect -10772 -394 -10770 -295
rect -10718 -394 -10716 -295
rect -10772 -567 -10716 -394
rect -10772 -700 -10716 -619
rect -10614 691 -10558 700
rect -10614 -394 -10612 385
rect -10560 -394 -10558 385
rect -10614 -700 -10558 -394
rect -10456 619 -10400 700
rect -10456 394 -10400 567
rect -10456 295 -10454 394
rect -10402 295 -10400 394
rect -10456 -394 -10454 -295
rect -10402 -394 -10400 -295
rect -10456 -567 -10400 -394
rect -10456 -700 -10400 -619
rect -10298 394 -10242 700
rect -10298 -385 -10296 394
rect -10244 -385 -10242 394
rect -10298 -700 -10242 -691
rect -10140 619 -10084 700
rect -10140 394 -10084 567
rect -10140 295 -10138 394
rect -10086 295 -10084 394
rect -10140 -394 -10138 -295
rect -10086 -394 -10084 -295
rect -10140 -567 -10084 -394
rect -10140 -700 -10084 -619
rect -9982 691 -9926 700
rect -9982 -394 -9980 385
rect -9928 -394 -9926 385
rect -9982 -700 -9926 -394
rect -9824 619 -9768 700
rect -9824 394 -9768 567
rect -9824 295 -9822 394
rect -9770 295 -9768 394
rect -9824 -394 -9822 -295
rect -9770 -394 -9768 -295
rect -9824 -567 -9768 -394
rect -9824 -700 -9768 -619
rect -9666 394 -9610 700
rect -9666 -385 -9664 394
rect -9612 -385 -9610 394
rect -9666 -700 -9610 -691
rect -9508 619 -9452 700
rect -9508 394 -9452 567
rect -9508 295 -9506 394
rect -9454 295 -9452 394
rect -9508 -394 -9506 -295
rect -9454 -394 -9452 -295
rect -9508 -567 -9452 -394
rect -9508 -700 -9452 -619
rect -9350 691 -9294 700
rect -9350 -394 -9348 385
rect -9296 -394 -9294 385
rect -9350 -700 -9294 -394
rect -9192 619 -9136 700
rect -9192 394 -9136 567
rect -9192 295 -9190 394
rect -9138 295 -9136 394
rect -9192 -394 -9190 -295
rect -9138 -394 -9136 -295
rect -9192 -567 -9136 -394
rect -9192 -700 -9136 -619
rect -9034 394 -8978 700
rect -9034 -385 -9032 394
rect -8980 -385 -8978 394
rect -9034 -700 -8978 -691
rect -8876 619 -8820 700
rect -8876 394 -8820 567
rect -8876 295 -8874 394
rect -8822 295 -8820 394
rect -8876 -394 -8874 -295
rect -8822 -394 -8820 -295
rect -8876 -567 -8820 -394
rect -8876 -700 -8820 -619
rect -8718 691 -8662 700
rect -8718 -394 -8716 385
rect -8664 -394 -8662 385
rect -8718 -700 -8662 -394
rect -8560 619 -8504 700
rect -8560 394 -8504 567
rect -8560 295 -8558 394
rect -8506 295 -8504 394
rect -8560 -394 -8558 -295
rect -8506 -394 -8504 -295
rect -8560 -567 -8504 -394
rect -8560 -700 -8504 -619
rect -8402 394 -8346 700
rect -8402 -385 -8400 394
rect -8348 -385 -8346 394
rect -8402 -700 -8346 -691
rect -8244 619 -8188 700
rect -8244 394 -8188 567
rect -8244 295 -8242 394
rect -8190 295 -8188 394
rect -8244 -394 -8242 -295
rect -8190 -394 -8188 -295
rect -8244 -567 -8188 -394
rect -8244 -700 -8188 -619
rect -8086 691 -8030 700
rect -8086 -394 -8084 385
rect -8032 -394 -8030 385
rect -8086 -700 -8030 -394
rect -7928 619 -7872 700
rect -7928 394 -7872 567
rect -7928 295 -7926 394
rect -7874 295 -7872 394
rect -7928 -394 -7926 -295
rect -7874 -394 -7872 -295
rect -7928 -567 -7872 -394
rect -7928 -700 -7872 -619
rect -7770 394 -7714 700
rect -7770 -385 -7768 394
rect -7716 -385 -7714 394
rect -7770 -700 -7714 -691
rect -7612 619 -7556 700
rect -7612 394 -7556 567
rect -7612 295 -7610 394
rect -7558 295 -7556 394
rect -7612 -394 -7610 -295
rect -7558 -394 -7556 -295
rect -7612 -567 -7556 -394
rect -7612 -700 -7556 -619
rect -7454 691 -7398 700
rect -7454 -394 -7452 385
rect -7400 -394 -7398 385
rect -7454 -700 -7398 -394
rect -7296 619 -7240 700
rect -7296 394 -7240 567
rect -7296 295 -7294 394
rect -7242 295 -7240 394
rect -7296 -394 -7294 -295
rect -7242 -394 -7240 -295
rect -7296 -567 -7240 -394
rect -7296 -700 -7240 -619
rect -7138 394 -7082 700
rect -7138 -385 -7136 394
rect -7084 -385 -7082 394
rect -7138 -700 -7082 -691
rect -6980 619 -6924 700
rect -6980 394 -6924 567
rect -6980 295 -6978 394
rect -6926 295 -6924 394
rect -6980 -394 -6978 -295
rect -6926 -394 -6924 -295
rect -6980 -567 -6924 -394
rect -6980 -700 -6924 -619
rect -6822 691 -6766 700
rect -6822 -394 -6820 385
rect -6768 -394 -6766 385
rect -6822 -700 -6766 -394
rect -6664 619 -6608 700
rect -6664 394 -6608 567
rect -6664 295 -6662 394
rect -6610 295 -6608 394
rect -6664 -394 -6662 -295
rect -6610 -394 -6608 -295
rect -6664 -567 -6608 -394
rect -6664 -700 -6608 -619
rect -6506 394 -6450 700
rect -6506 -385 -6504 394
rect -6452 -385 -6450 394
rect -6506 -700 -6450 -691
rect -6348 619 -6292 700
rect -6348 394 -6292 567
rect -6348 295 -6346 394
rect -6294 295 -6292 394
rect -6348 -394 -6346 -295
rect -6294 -394 -6292 -295
rect -6348 -567 -6292 -394
rect -6348 -700 -6292 -619
rect -6190 691 -6134 700
rect -6190 -394 -6188 385
rect -6136 -394 -6134 385
rect -6190 -700 -6134 -394
rect -6032 619 -5976 700
rect -6032 394 -5976 567
rect -6032 295 -6030 394
rect -5978 295 -5976 394
rect -6032 -394 -6030 -295
rect -5978 -394 -5976 -295
rect -6032 -567 -5976 -394
rect -6032 -700 -5976 -619
rect -5874 394 -5818 700
rect -5874 -385 -5872 394
rect -5820 -385 -5818 394
rect -5874 -700 -5818 -691
rect -5716 619 -5660 700
rect -5716 394 -5660 567
rect -5716 295 -5714 394
rect -5662 295 -5660 394
rect -5716 -394 -5714 -295
rect -5662 -394 -5660 -295
rect -5716 -567 -5660 -394
rect -5716 -700 -5660 -619
rect -5558 691 -5502 700
rect -5558 -394 -5556 385
rect -5504 -394 -5502 385
rect -5558 -700 -5502 -394
rect -5400 619 -5344 700
rect -5400 394 -5344 567
rect -5400 295 -5398 394
rect -5346 295 -5344 394
rect -5400 -394 -5398 -295
rect -5346 -394 -5344 -295
rect -5400 -567 -5344 -394
rect -5400 -700 -5344 -619
rect -5242 394 -5186 700
rect -5242 -385 -5240 394
rect -5188 -385 -5186 394
rect -5242 -700 -5186 -691
rect -5084 619 -5028 700
rect -5084 394 -5028 567
rect -5084 295 -5082 394
rect -5030 295 -5028 394
rect -5084 -394 -5082 -295
rect -5030 -394 -5028 -295
rect -5084 -567 -5028 -394
rect -5084 -700 -5028 -619
rect -4926 691 -4870 700
rect -4926 -394 -4924 385
rect -4872 -394 -4870 385
rect -4926 -700 -4870 -394
rect -4768 619 -4712 700
rect -4768 394 -4712 567
rect -4768 295 -4766 394
rect -4714 295 -4712 394
rect -4768 -394 -4766 -295
rect -4714 -394 -4712 -295
rect -4768 -567 -4712 -394
rect -4768 -700 -4712 -619
rect -4452 619 -4396 700
rect -4452 394 -4396 567
rect -4452 295 -4450 394
rect -4398 295 -4396 394
rect -4452 -394 -4450 -295
rect -4398 -394 -4396 -295
rect -4452 -567 -4396 -394
rect -4452 -700 -4396 -619
rect -4294 394 -4238 700
rect -4294 -385 -4292 394
rect -4240 -385 -4238 394
rect -4294 -700 -4238 -691
rect -4136 619 -4080 700
rect -4136 394 -4080 567
rect -4136 295 -4134 394
rect -4082 295 -4080 394
rect -4136 -394 -4134 -295
rect -4082 -394 -4080 -295
rect -4136 -567 -4080 -394
rect -4136 -700 -4080 -619
rect -3978 691 -3922 700
rect -3978 -394 -3976 385
rect -3924 -394 -3922 385
rect -3978 -700 -3922 -394
rect -3820 619 -3764 700
rect -3820 394 -3764 567
rect -3820 295 -3818 394
rect -3766 295 -3764 394
rect -3820 -394 -3818 -295
rect -3766 -394 -3764 -295
rect -3820 -567 -3764 -394
rect -3820 -700 -3764 -619
rect -3662 394 -3606 700
rect -3662 -385 -3660 394
rect -3608 -385 -3606 394
rect -3662 -700 -3606 -691
rect -3504 619 -3448 700
rect -3504 394 -3448 567
rect -3504 295 -3502 394
rect -3450 295 -3448 394
rect -3504 -394 -3502 -295
rect -3450 -394 -3448 -295
rect -3504 -567 -3448 -394
rect -3504 -700 -3448 -619
rect -3346 691 -3290 700
rect -3346 -394 -3344 385
rect -3292 -394 -3290 385
rect -3346 -700 -3290 -394
rect -3188 619 -3132 700
rect -3188 394 -3132 567
rect -3188 295 -3186 394
rect -3134 295 -3132 394
rect -3188 -394 -3186 -295
rect -3134 -394 -3132 -295
rect -3188 -567 -3132 -394
rect -3188 -700 -3132 -619
rect -3030 394 -2974 700
rect -3030 -385 -3028 394
rect -2976 -385 -2974 394
rect -3030 -700 -2974 -691
rect -2872 619 -2816 700
rect -2872 394 -2816 567
rect -2872 295 -2870 394
rect -2818 295 -2816 394
rect -2872 -394 -2870 -295
rect -2818 -394 -2816 -295
rect -2872 -567 -2816 -394
rect -2872 -700 -2816 -619
rect -2714 691 -2658 700
rect -2714 -394 -2712 385
rect -2660 -394 -2658 385
rect -2714 -700 -2658 -394
rect -2556 619 -2500 700
rect -2556 394 -2500 567
rect -2556 295 -2554 394
rect -2502 295 -2500 394
rect -2556 -394 -2554 -295
rect -2502 -394 -2500 -295
rect -2556 -567 -2500 -394
rect -2556 -700 -2500 -619
rect -2398 394 -2342 700
rect -2398 -385 -2396 394
rect -2344 -385 -2342 394
rect -2398 -700 -2342 -691
rect -2240 619 -2184 700
rect -2240 394 -2184 567
rect -2240 295 -2238 394
rect -2186 295 -2184 394
rect -2240 -394 -2238 -295
rect -2186 -394 -2184 -295
rect -2240 -567 -2184 -394
rect -2240 -700 -2184 -619
rect -2082 691 -2026 700
rect -2082 -394 -2080 385
rect -2028 -394 -2026 385
rect -2082 -700 -2026 -394
rect -1924 619 -1868 700
rect -1924 394 -1868 567
rect -1924 295 -1922 394
rect -1870 295 -1868 394
rect -1924 -394 -1922 -295
rect -1870 -394 -1868 -295
rect -1924 -567 -1868 -394
rect -1924 -700 -1868 -619
rect -1766 394 -1710 700
rect -1766 -385 -1764 394
rect -1712 -385 -1710 394
rect -1766 -700 -1710 -691
rect -1608 619 -1552 700
rect -1608 394 -1552 567
rect -1608 295 -1606 394
rect -1554 295 -1552 394
rect -1608 -394 -1606 -295
rect -1554 -394 -1552 -295
rect -1608 -567 -1552 -394
rect -1608 -700 -1552 -619
rect -1450 691 -1394 700
rect -1450 -394 -1448 385
rect -1396 -394 -1394 385
rect -1450 -700 -1394 -394
rect -1292 619 -1236 700
rect -1292 394 -1236 567
rect -1292 295 -1290 394
rect -1238 295 -1236 394
rect -1292 -394 -1290 -295
rect -1238 -394 -1236 -295
rect -1292 -567 -1236 -394
rect -1292 -700 -1236 -619
rect -1134 394 -1078 700
rect -1134 -385 -1132 394
rect -1080 -385 -1078 394
rect -1134 -700 -1078 -691
rect -976 619 -920 700
rect -976 394 -920 567
rect -976 295 -974 394
rect -922 295 -920 394
rect -976 -394 -974 -295
rect -922 -394 -920 -295
rect -976 -567 -920 -394
rect -976 -700 -920 -619
rect -818 691 -762 700
rect -818 -394 -816 385
rect -764 -394 -762 385
rect -818 -700 -762 -394
rect -660 619 -604 700
rect -660 394 -604 567
rect -660 295 -658 394
rect -606 295 -604 394
rect -660 -394 -658 -295
rect -606 -394 -604 -295
rect -660 -567 -604 -394
rect -660 -700 -604 -619
rect -502 394 -446 700
rect -502 -385 -500 394
rect -448 -385 -446 394
rect -502 -700 -446 -691
rect -344 619 -288 700
rect -344 394 -288 567
rect -344 295 -342 394
rect -290 295 -288 394
rect -344 -394 -342 -295
rect -290 -394 -288 -295
rect -344 -567 -288 -394
rect -344 -700 -288 -619
rect -186 691 -130 700
rect -186 -394 -184 385
rect -132 -394 -130 385
rect -186 -700 -130 -394
rect -28 619 28 700
rect -28 394 28 567
rect -28 295 -26 394
rect 26 295 28 394
rect -28 -394 -26 -295
rect 26 -394 28 -295
rect -28 -567 28 -394
rect -28 -700 28 -619
rect 130 691 186 700
rect 130 -394 132 385
rect 184 -394 186 385
rect 130 -700 186 -394
rect 288 619 344 700
rect 288 394 344 567
rect 288 295 290 394
rect 342 295 344 394
rect 288 -394 290 -295
rect 342 -394 344 -295
rect 288 -567 344 -394
rect 288 -700 344 -619
rect 446 394 502 700
rect 446 -385 448 394
rect 500 -385 502 394
rect 446 -700 502 -691
rect 604 619 660 700
rect 604 394 660 567
rect 604 295 606 394
rect 658 295 660 394
rect 604 -394 606 -295
rect 658 -394 660 -295
rect 604 -567 660 -394
rect 604 -700 660 -619
rect 762 691 818 700
rect 762 -394 764 385
rect 816 -394 818 385
rect 762 -700 818 -394
rect 920 619 976 700
rect 920 394 976 567
rect 920 295 922 394
rect 974 295 976 394
rect 920 -394 922 -295
rect 974 -394 976 -295
rect 920 -567 976 -394
rect 920 -700 976 -619
rect 1078 394 1134 700
rect 1078 -385 1080 394
rect 1132 -385 1134 394
rect 1078 -700 1134 -691
rect 1236 619 1292 700
rect 1236 394 1292 567
rect 1236 295 1238 394
rect 1290 295 1292 394
rect 1236 -394 1238 -295
rect 1290 -394 1292 -295
rect 1236 -567 1292 -394
rect 1236 -700 1292 -619
rect 1394 691 1450 700
rect 1394 -394 1396 385
rect 1448 -394 1450 385
rect 1394 -700 1450 -394
rect 1552 619 1608 700
rect 1552 394 1608 567
rect 1552 295 1554 394
rect 1606 295 1608 394
rect 1552 -394 1554 -295
rect 1606 -394 1608 -295
rect 1552 -567 1608 -394
rect 1552 -700 1608 -619
rect 1710 394 1766 700
rect 1710 -385 1712 394
rect 1764 -385 1766 394
rect 1710 -700 1766 -691
rect 1868 619 1924 700
rect 1868 394 1924 567
rect 1868 295 1870 394
rect 1922 295 1924 394
rect 1868 -394 1870 -295
rect 1922 -394 1924 -295
rect 1868 -567 1924 -394
rect 1868 -700 1924 -619
rect 2026 691 2082 700
rect 2026 -394 2028 385
rect 2080 -394 2082 385
rect 2026 -700 2082 -394
rect 2184 619 2240 700
rect 2184 394 2240 567
rect 2184 295 2186 394
rect 2238 295 2240 394
rect 2184 -394 2186 -295
rect 2238 -394 2240 -295
rect 2184 -567 2240 -394
rect 2184 -700 2240 -619
rect 2342 394 2398 700
rect 2342 -385 2344 394
rect 2396 -385 2398 394
rect 2342 -700 2398 -691
rect 2500 619 2556 700
rect 2500 394 2556 567
rect 2500 295 2502 394
rect 2554 295 2556 394
rect 2500 -394 2502 -295
rect 2554 -394 2556 -295
rect 2500 -567 2556 -394
rect 2500 -700 2556 -619
rect 2658 691 2714 700
rect 2658 -394 2660 385
rect 2712 -394 2714 385
rect 2658 -700 2714 -394
rect 2816 619 2872 700
rect 2816 394 2872 567
rect 2816 295 2818 394
rect 2870 295 2872 394
rect 2816 -394 2818 -295
rect 2870 -394 2872 -295
rect 2816 -567 2872 -394
rect 2816 -700 2872 -619
rect 2974 394 3030 700
rect 2974 -385 2976 394
rect 3028 -385 3030 394
rect 2974 -700 3030 -691
rect 3132 619 3188 700
rect 3132 394 3188 567
rect 3132 295 3134 394
rect 3186 295 3188 394
rect 3132 -394 3134 -295
rect 3186 -394 3188 -295
rect 3132 -567 3188 -394
rect 3132 -700 3188 -619
rect 3290 691 3346 700
rect 3290 -394 3292 385
rect 3344 -394 3346 385
rect 3290 -700 3346 -394
rect 3448 619 3504 700
rect 3448 394 3504 567
rect 3448 295 3450 394
rect 3502 295 3504 394
rect 3448 -394 3450 -295
rect 3502 -394 3504 -295
rect 3448 -567 3504 -394
rect 3448 -700 3504 -619
rect 3606 394 3662 700
rect 3606 -385 3608 394
rect 3660 -385 3662 394
rect 3606 -700 3662 -691
rect 3764 619 3820 700
rect 3764 394 3820 567
rect 3764 295 3766 394
rect 3818 295 3820 394
rect 3764 -394 3766 -295
rect 3818 -394 3820 -295
rect 3764 -567 3820 -394
rect 3764 -700 3820 -619
rect 3922 691 3978 700
rect 3922 -394 3924 385
rect 3976 -394 3978 385
rect 3922 -700 3978 -394
rect 4080 619 4136 700
rect 4080 394 4136 567
rect 4080 295 4082 394
rect 4134 295 4136 394
rect 4080 -394 4082 -295
rect 4134 -394 4136 -295
rect 4080 -567 4136 -394
rect 4080 -700 4136 -619
rect 4238 394 4294 700
rect 4238 -385 4240 394
rect 4292 -385 4294 394
rect 4238 -700 4294 -691
rect 4396 619 4452 700
rect 4396 394 4452 567
rect 4396 295 4398 394
rect 4450 295 4452 394
rect 4396 -394 4398 -295
rect 4450 -394 4452 -295
rect 4396 -567 4452 -394
rect 4396 -700 4452 -619
rect 4712 619 4768 700
rect 4712 394 4768 567
rect 4712 295 4714 394
rect 4766 295 4768 394
rect 4712 -394 4714 -295
rect 4766 -394 4768 -295
rect 4712 -567 4768 -394
rect 4712 -700 4768 -619
rect 4870 691 4926 700
rect 4870 -394 4872 385
rect 4924 -394 4926 385
rect 4870 -700 4926 -394
rect 5028 619 5084 700
rect 5028 394 5084 567
rect 5028 295 5030 394
rect 5082 295 5084 394
rect 5028 -394 5030 -295
rect 5082 -394 5084 -295
rect 5028 -567 5084 -394
rect 5028 -700 5084 -619
rect 5186 394 5242 700
rect 5186 -385 5188 394
rect 5240 -385 5242 394
rect 5186 -700 5242 -691
rect 5344 619 5400 700
rect 5344 394 5400 567
rect 5344 295 5346 394
rect 5398 295 5400 394
rect 5344 -394 5346 -295
rect 5398 -394 5400 -295
rect 5344 -567 5400 -394
rect 5344 -700 5400 -619
rect 5502 691 5558 700
rect 5502 -394 5504 385
rect 5556 -394 5558 385
rect 5502 -700 5558 -394
rect 5660 619 5716 700
rect 5660 394 5716 567
rect 5660 295 5662 394
rect 5714 295 5716 394
rect 5660 -394 5662 -295
rect 5714 -394 5716 -295
rect 5660 -567 5716 -394
rect 5660 -700 5716 -619
rect 5818 394 5874 700
rect 5818 -385 5820 394
rect 5872 -385 5874 394
rect 5818 -700 5874 -691
rect 5976 619 6032 700
rect 5976 394 6032 567
rect 5976 295 5978 394
rect 6030 295 6032 394
rect 5976 -394 5978 -295
rect 6030 -394 6032 -295
rect 5976 -567 6032 -394
rect 5976 -700 6032 -619
rect 6134 691 6190 700
rect 6134 -394 6136 385
rect 6188 -394 6190 385
rect 6134 -700 6190 -394
rect 6292 619 6348 700
rect 6292 394 6348 567
rect 6292 295 6294 394
rect 6346 295 6348 394
rect 6292 -394 6294 -295
rect 6346 -394 6348 -295
rect 6292 -567 6348 -394
rect 6292 -700 6348 -619
rect 6450 394 6506 700
rect 6450 -385 6452 394
rect 6504 -385 6506 394
rect 6450 -700 6506 -691
rect 6608 619 6664 700
rect 6608 394 6664 567
rect 6608 295 6610 394
rect 6662 295 6664 394
rect 6608 -394 6610 -295
rect 6662 -394 6664 -295
rect 6608 -567 6664 -394
rect 6608 -700 6664 -619
rect 6766 691 6822 700
rect 6766 -394 6768 385
rect 6820 -394 6822 385
rect 6766 -700 6822 -394
rect 6924 619 6980 700
rect 6924 394 6980 567
rect 6924 295 6926 394
rect 6978 295 6980 394
rect 6924 -394 6926 -295
rect 6978 -394 6980 -295
rect 6924 -567 6980 -394
rect 6924 -700 6980 -619
rect 7082 394 7138 700
rect 7082 -385 7084 394
rect 7136 -385 7138 394
rect 7082 -700 7138 -691
rect 7240 619 7296 700
rect 7240 394 7296 567
rect 7240 295 7242 394
rect 7294 295 7296 394
rect 7240 -394 7242 -295
rect 7294 -394 7296 -295
rect 7240 -567 7296 -394
rect 7240 -700 7296 -619
rect 7398 691 7454 700
rect 7398 -394 7400 385
rect 7452 -394 7454 385
rect 7398 -700 7454 -394
rect 7556 619 7612 700
rect 7556 394 7612 567
rect 7556 295 7558 394
rect 7610 295 7612 394
rect 7556 -394 7558 -295
rect 7610 -394 7612 -295
rect 7556 -567 7612 -394
rect 7556 -700 7612 -619
rect 7714 394 7770 700
rect 7714 -385 7716 394
rect 7768 -385 7770 394
rect 7714 -700 7770 -691
rect 7872 619 7928 700
rect 7872 394 7928 567
rect 7872 295 7874 394
rect 7926 295 7928 394
rect 7872 -394 7874 -295
rect 7926 -394 7928 -295
rect 7872 -567 7928 -394
rect 7872 -700 7928 -619
rect 8030 691 8086 700
rect 8030 -394 8032 385
rect 8084 -394 8086 385
rect 8030 -700 8086 -394
rect 8188 619 8244 700
rect 8188 394 8244 567
rect 8188 295 8190 394
rect 8242 295 8244 394
rect 8188 -394 8190 -295
rect 8242 -394 8244 -295
rect 8188 -567 8244 -394
rect 8188 -700 8244 -619
rect 8346 394 8402 700
rect 8346 -385 8348 394
rect 8400 -385 8402 394
rect 8346 -700 8402 -691
rect 8504 619 8560 700
rect 8504 394 8560 567
rect 8504 295 8506 394
rect 8558 295 8560 394
rect 8504 -394 8506 -295
rect 8558 -394 8560 -295
rect 8504 -567 8560 -394
rect 8504 -700 8560 -619
rect 8662 691 8718 700
rect 8662 -394 8664 385
rect 8716 -394 8718 385
rect 8662 -700 8718 -394
rect 8820 619 8876 700
rect 8820 394 8876 567
rect 8820 295 8822 394
rect 8874 295 8876 394
rect 8820 -394 8822 -295
rect 8874 -394 8876 -295
rect 8820 -567 8876 -394
rect 8820 -700 8876 -619
rect 8978 394 9034 700
rect 8978 -385 8980 394
rect 9032 -385 9034 394
rect 8978 -700 9034 -691
rect 9136 619 9192 700
rect 9136 394 9192 567
rect 9136 295 9138 394
rect 9190 295 9192 394
rect 9136 -394 9138 -295
rect 9190 -394 9192 -295
rect 9136 -567 9192 -394
rect 9136 -700 9192 -619
rect 9294 691 9350 700
rect 9294 -394 9296 385
rect 9348 -394 9350 385
rect 9294 -700 9350 -394
rect 9452 619 9508 700
rect 9452 394 9508 567
rect 9452 295 9454 394
rect 9506 295 9508 394
rect 9452 -394 9454 -295
rect 9506 -394 9508 -295
rect 9452 -567 9508 -394
rect 9452 -700 9508 -619
rect 9610 394 9666 700
rect 9610 -385 9612 394
rect 9664 -385 9666 394
rect 9610 -700 9666 -691
rect 9768 619 9824 700
rect 9768 394 9824 567
rect 9768 295 9770 394
rect 9822 295 9824 394
rect 9768 -394 9770 -295
rect 9822 -394 9824 -295
rect 9768 -567 9824 -394
rect 9768 -700 9824 -619
rect 9926 691 9982 700
rect 9926 -394 9928 385
rect 9980 -394 9982 385
rect 9926 -700 9982 -394
rect 10084 619 10140 700
rect 10084 394 10140 567
rect 10084 295 10086 394
rect 10138 295 10140 394
rect 10084 -394 10086 -295
rect 10138 -394 10140 -295
rect 10084 -567 10140 -394
rect 10084 -700 10140 -619
rect 10242 394 10298 700
rect 10242 -385 10244 394
rect 10296 -385 10298 394
rect 10242 -700 10298 -691
rect 10400 619 10456 700
rect 10400 394 10456 567
rect 10400 295 10402 394
rect 10454 295 10456 394
rect 10400 -394 10402 -295
rect 10454 -394 10456 -295
rect 10400 -567 10456 -394
rect 10400 -700 10456 -619
rect 10558 691 10614 700
rect 10558 -394 10560 385
rect 10612 -394 10614 385
rect 10558 -700 10614 -394
rect 10716 619 10772 700
rect 10716 394 10772 567
rect 10716 295 10718 394
rect 10770 295 10772 394
rect 10716 -394 10718 -295
rect 10770 -394 10772 -295
rect 10716 -567 10772 -394
rect 10716 -700 10772 -619
rect 10874 394 10930 700
rect 10874 -385 10876 394
rect 10928 -385 10930 394
rect 10874 -700 10930 -691
rect 11032 619 11088 700
rect 11032 394 11088 567
rect 11032 295 11034 394
rect 11086 295 11088 394
rect 11032 -394 11034 -295
rect 11086 -394 11088 -295
rect 11032 -567 11088 -394
rect 11032 -700 11088 -619
rect 11190 691 11246 700
rect 11190 -394 11192 385
rect 11244 -394 11246 385
rect 11190 -700 11246 -394
rect 11348 619 11404 700
rect 11348 394 11404 567
rect 11348 295 11350 394
rect 11402 295 11404 394
rect 11348 -394 11350 -295
rect 11402 -394 11404 -295
rect 11348 -567 11404 -394
rect 11348 -700 11404 -619
rect 11506 394 11562 700
rect 11506 -385 11508 394
rect 11560 -385 11562 394
rect 11506 -700 11562 -691
rect 11664 619 11720 700
rect 11664 394 11720 567
rect 11664 295 11666 394
rect 11718 295 11720 394
rect 11664 -394 11666 -295
rect 11718 -394 11720 -295
rect 11664 -567 11720 -394
rect 11664 -700 11720 -619
rect 11822 691 11878 700
rect 11822 -394 11824 385
rect 11876 -394 11878 385
rect 11822 -700 11878 -394
rect 11980 619 12036 700
rect 11980 394 12036 567
rect 11980 295 11982 394
rect 12034 295 12036 394
rect 11980 -394 11982 -295
rect 12034 -394 12036 -295
rect 11980 -567 12036 -394
rect 11980 -700 12036 -619
rect 12138 394 12194 700
rect 12138 -385 12140 394
rect 12192 -385 12194 394
rect 12138 -700 12194 -691
rect 12296 619 12352 700
rect 12296 394 12352 567
rect 12296 295 12298 394
rect 12350 295 12352 394
rect 12296 -394 12298 -295
rect 12350 -394 12352 -295
rect 12296 -567 12352 -394
rect 12296 -700 12352 -619
rect 12454 691 12510 700
rect 12454 -394 12456 385
rect 12508 -394 12510 385
rect 12454 -700 12510 -394
rect 12612 619 12668 700
rect 12612 394 12668 567
rect 12612 295 12614 394
rect 12666 295 12668 394
rect 12612 -394 12614 -295
rect 12666 -394 12668 -295
rect 12612 -567 12668 -394
rect 12612 -700 12668 -619
rect 12770 394 12826 700
rect 12770 -385 12772 394
rect 12824 -385 12826 394
rect 12770 -700 12826 -691
rect 12928 619 12984 700
rect 12928 394 12984 567
rect 12928 295 12930 394
rect 12982 295 12984 394
rect 12928 -394 12930 -295
rect 12982 -394 12984 -295
rect 12928 -567 12984 -394
rect 12928 -700 12984 -619
<< via2 >>
rect -12984 -295 -12982 295
rect -12982 -295 -12930 295
rect -12930 -295 -12928 295
rect -12826 -394 -12824 -385
rect -12824 -394 -12772 -385
rect -12772 -394 -12770 -385
rect -12826 -691 -12770 -394
rect -12668 -295 -12666 295
rect -12666 -295 -12614 295
rect -12614 -295 -12612 295
rect -12510 394 -12454 691
rect -12510 385 -12508 394
rect -12508 385 -12456 394
rect -12456 385 -12454 394
rect -12352 -295 -12350 295
rect -12350 -295 -12298 295
rect -12298 -295 -12296 295
rect -12194 -394 -12192 -385
rect -12192 -394 -12140 -385
rect -12140 -394 -12138 -385
rect -12194 -691 -12138 -394
rect -12036 -295 -12034 295
rect -12034 -295 -11982 295
rect -11982 -295 -11980 295
rect -11878 394 -11822 691
rect -11878 385 -11876 394
rect -11876 385 -11824 394
rect -11824 385 -11822 394
rect -11720 -295 -11718 295
rect -11718 -295 -11666 295
rect -11666 -295 -11664 295
rect -11562 -394 -11560 -385
rect -11560 -394 -11508 -385
rect -11508 -394 -11506 -385
rect -11562 -691 -11506 -394
rect -11404 -295 -11402 295
rect -11402 -295 -11350 295
rect -11350 -295 -11348 295
rect -11246 394 -11190 691
rect -11246 385 -11244 394
rect -11244 385 -11192 394
rect -11192 385 -11190 394
rect -11088 -295 -11086 295
rect -11086 -295 -11034 295
rect -11034 -295 -11032 295
rect -10930 -394 -10928 -385
rect -10928 -394 -10876 -385
rect -10876 -394 -10874 -385
rect -10930 -691 -10874 -394
rect -10772 -295 -10770 295
rect -10770 -295 -10718 295
rect -10718 -295 -10716 295
rect -10614 394 -10558 691
rect -10614 385 -10612 394
rect -10612 385 -10560 394
rect -10560 385 -10558 394
rect -10456 -295 -10454 295
rect -10454 -295 -10402 295
rect -10402 -295 -10400 295
rect -10298 -394 -10296 -385
rect -10296 -394 -10244 -385
rect -10244 -394 -10242 -385
rect -10298 -691 -10242 -394
rect -10140 -295 -10138 295
rect -10138 -295 -10086 295
rect -10086 -295 -10084 295
rect -9982 394 -9926 691
rect -9982 385 -9980 394
rect -9980 385 -9928 394
rect -9928 385 -9926 394
rect -9824 -295 -9822 295
rect -9822 -295 -9770 295
rect -9770 -295 -9768 295
rect -9666 -394 -9664 -385
rect -9664 -394 -9612 -385
rect -9612 -394 -9610 -385
rect -9666 -691 -9610 -394
rect -9508 -295 -9506 295
rect -9506 -295 -9454 295
rect -9454 -295 -9452 295
rect -9350 394 -9294 691
rect -9350 385 -9348 394
rect -9348 385 -9296 394
rect -9296 385 -9294 394
rect -9192 -295 -9190 295
rect -9190 -295 -9138 295
rect -9138 -295 -9136 295
rect -9034 -394 -9032 -385
rect -9032 -394 -8980 -385
rect -8980 -394 -8978 -385
rect -9034 -691 -8978 -394
rect -8876 -295 -8874 295
rect -8874 -295 -8822 295
rect -8822 -295 -8820 295
rect -8718 394 -8662 691
rect -8718 385 -8716 394
rect -8716 385 -8664 394
rect -8664 385 -8662 394
rect -8560 -295 -8558 295
rect -8558 -295 -8506 295
rect -8506 -295 -8504 295
rect -8402 -394 -8400 -385
rect -8400 -394 -8348 -385
rect -8348 -394 -8346 -385
rect -8402 -691 -8346 -394
rect -8244 -295 -8242 295
rect -8242 -295 -8190 295
rect -8190 -295 -8188 295
rect -8086 394 -8030 691
rect -8086 385 -8084 394
rect -8084 385 -8032 394
rect -8032 385 -8030 394
rect -7928 -295 -7926 295
rect -7926 -295 -7874 295
rect -7874 -295 -7872 295
rect -7770 -394 -7768 -385
rect -7768 -394 -7716 -385
rect -7716 -394 -7714 -385
rect -7770 -691 -7714 -394
rect -7612 -295 -7610 295
rect -7610 -295 -7558 295
rect -7558 -295 -7556 295
rect -7454 394 -7398 691
rect -7454 385 -7452 394
rect -7452 385 -7400 394
rect -7400 385 -7398 394
rect -7296 -295 -7294 295
rect -7294 -295 -7242 295
rect -7242 -295 -7240 295
rect -7138 -394 -7136 -385
rect -7136 -394 -7084 -385
rect -7084 -394 -7082 -385
rect -7138 -691 -7082 -394
rect -6980 -295 -6978 295
rect -6978 -295 -6926 295
rect -6926 -295 -6924 295
rect -6822 394 -6766 691
rect -6822 385 -6820 394
rect -6820 385 -6768 394
rect -6768 385 -6766 394
rect -6664 -295 -6662 295
rect -6662 -295 -6610 295
rect -6610 -295 -6608 295
rect -6506 -394 -6504 -385
rect -6504 -394 -6452 -385
rect -6452 -394 -6450 -385
rect -6506 -691 -6450 -394
rect -6348 -295 -6346 295
rect -6346 -295 -6294 295
rect -6294 -295 -6292 295
rect -6190 394 -6134 691
rect -6190 385 -6188 394
rect -6188 385 -6136 394
rect -6136 385 -6134 394
rect -6032 -295 -6030 295
rect -6030 -295 -5978 295
rect -5978 -295 -5976 295
rect -5874 -394 -5872 -385
rect -5872 -394 -5820 -385
rect -5820 -394 -5818 -385
rect -5874 -691 -5818 -394
rect -5716 -295 -5714 295
rect -5714 -295 -5662 295
rect -5662 -295 -5660 295
rect -5558 394 -5502 691
rect -5558 385 -5556 394
rect -5556 385 -5504 394
rect -5504 385 -5502 394
rect -5400 -295 -5398 295
rect -5398 -295 -5346 295
rect -5346 -295 -5344 295
rect -5242 -394 -5240 -385
rect -5240 -394 -5188 -385
rect -5188 -394 -5186 -385
rect -5242 -691 -5186 -394
rect -5084 -295 -5082 295
rect -5082 -295 -5030 295
rect -5030 -295 -5028 295
rect -4926 394 -4870 691
rect -4926 385 -4924 394
rect -4924 385 -4872 394
rect -4872 385 -4870 394
rect -4768 -295 -4766 295
rect -4766 -295 -4714 295
rect -4714 -295 -4712 295
rect -4452 -295 -4450 295
rect -4450 -295 -4398 295
rect -4398 -295 -4396 295
rect -4294 -394 -4292 -385
rect -4292 -394 -4240 -385
rect -4240 -394 -4238 -385
rect -4294 -691 -4238 -394
rect -4136 -295 -4134 295
rect -4134 -295 -4082 295
rect -4082 -295 -4080 295
rect -3978 394 -3922 691
rect -3978 385 -3976 394
rect -3976 385 -3924 394
rect -3924 385 -3922 394
rect -3820 -295 -3818 295
rect -3818 -295 -3766 295
rect -3766 -295 -3764 295
rect -3662 -394 -3660 -385
rect -3660 -394 -3608 -385
rect -3608 -394 -3606 -385
rect -3662 -691 -3606 -394
rect -3504 -295 -3502 295
rect -3502 -295 -3450 295
rect -3450 -295 -3448 295
rect -3346 394 -3290 691
rect -3346 385 -3344 394
rect -3344 385 -3292 394
rect -3292 385 -3290 394
rect -3188 -295 -3186 295
rect -3186 -295 -3134 295
rect -3134 -295 -3132 295
rect -3030 -394 -3028 -385
rect -3028 -394 -2976 -385
rect -2976 -394 -2974 -385
rect -3030 -691 -2974 -394
rect -2872 -295 -2870 295
rect -2870 -295 -2818 295
rect -2818 -295 -2816 295
rect -2714 394 -2658 691
rect -2714 385 -2712 394
rect -2712 385 -2660 394
rect -2660 385 -2658 394
rect -2556 -295 -2554 295
rect -2554 -295 -2502 295
rect -2502 -295 -2500 295
rect -2398 -394 -2396 -385
rect -2396 -394 -2344 -385
rect -2344 -394 -2342 -385
rect -2398 -691 -2342 -394
rect -2240 -295 -2238 295
rect -2238 -295 -2186 295
rect -2186 -295 -2184 295
rect -2082 394 -2026 691
rect -2082 385 -2080 394
rect -2080 385 -2028 394
rect -2028 385 -2026 394
rect -1924 -295 -1922 295
rect -1922 -295 -1870 295
rect -1870 -295 -1868 295
rect -1766 -394 -1764 -385
rect -1764 -394 -1712 -385
rect -1712 -394 -1710 -385
rect -1766 -691 -1710 -394
rect -1608 -295 -1606 295
rect -1606 -295 -1554 295
rect -1554 -295 -1552 295
rect -1450 394 -1394 691
rect -1450 385 -1448 394
rect -1448 385 -1396 394
rect -1396 385 -1394 394
rect -1292 -295 -1290 295
rect -1290 -295 -1238 295
rect -1238 -295 -1236 295
rect -1134 -394 -1132 -385
rect -1132 -394 -1080 -385
rect -1080 -394 -1078 -385
rect -1134 -691 -1078 -394
rect -976 -295 -974 295
rect -974 -295 -922 295
rect -922 -295 -920 295
rect -818 394 -762 691
rect -818 385 -816 394
rect -816 385 -764 394
rect -764 385 -762 394
rect -660 -295 -658 295
rect -658 -295 -606 295
rect -606 -295 -604 295
rect -502 -394 -500 -385
rect -500 -394 -448 -385
rect -448 -394 -446 -385
rect -502 -691 -446 -394
rect -344 -295 -342 295
rect -342 -295 -290 295
rect -290 -295 -288 295
rect -186 394 -130 691
rect -186 385 -184 394
rect -184 385 -132 394
rect -132 385 -130 394
rect -28 -295 -26 295
rect -26 -295 26 295
rect 26 -295 28 295
rect 130 394 186 691
rect 130 385 132 394
rect 132 385 184 394
rect 184 385 186 394
rect 288 -295 290 295
rect 290 -295 342 295
rect 342 -295 344 295
rect 446 -394 448 -385
rect 448 -394 500 -385
rect 500 -394 502 -385
rect 446 -691 502 -394
rect 604 -295 606 295
rect 606 -295 658 295
rect 658 -295 660 295
rect 762 394 818 691
rect 762 385 764 394
rect 764 385 816 394
rect 816 385 818 394
rect 920 -295 922 295
rect 922 -295 974 295
rect 974 -295 976 295
rect 1078 -394 1080 -385
rect 1080 -394 1132 -385
rect 1132 -394 1134 -385
rect 1078 -691 1134 -394
rect 1236 -295 1238 295
rect 1238 -295 1290 295
rect 1290 -295 1292 295
rect 1394 394 1450 691
rect 1394 385 1396 394
rect 1396 385 1448 394
rect 1448 385 1450 394
rect 1552 -295 1554 295
rect 1554 -295 1606 295
rect 1606 -295 1608 295
rect 1710 -394 1712 -385
rect 1712 -394 1764 -385
rect 1764 -394 1766 -385
rect 1710 -691 1766 -394
rect 1868 -295 1870 295
rect 1870 -295 1922 295
rect 1922 -295 1924 295
rect 2026 394 2082 691
rect 2026 385 2028 394
rect 2028 385 2080 394
rect 2080 385 2082 394
rect 2184 -295 2186 295
rect 2186 -295 2238 295
rect 2238 -295 2240 295
rect 2342 -394 2344 -385
rect 2344 -394 2396 -385
rect 2396 -394 2398 -385
rect 2342 -691 2398 -394
rect 2500 -295 2502 295
rect 2502 -295 2554 295
rect 2554 -295 2556 295
rect 2658 394 2714 691
rect 2658 385 2660 394
rect 2660 385 2712 394
rect 2712 385 2714 394
rect 2816 -295 2818 295
rect 2818 -295 2870 295
rect 2870 -295 2872 295
rect 2974 -394 2976 -385
rect 2976 -394 3028 -385
rect 3028 -394 3030 -385
rect 2974 -691 3030 -394
rect 3132 -295 3134 295
rect 3134 -295 3186 295
rect 3186 -295 3188 295
rect 3290 394 3346 691
rect 3290 385 3292 394
rect 3292 385 3344 394
rect 3344 385 3346 394
rect 3448 -295 3450 295
rect 3450 -295 3502 295
rect 3502 -295 3504 295
rect 3606 -394 3608 -385
rect 3608 -394 3660 -385
rect 3660 -394 3662 -385
rect 3606 -691 3662 -394
rect 3764 -295 3766 295
rect 3766 -295 3818 295
rect 3818 -295 3820 295
rect 3922 394 3978 691
rect 3922 385 3924 394
rect 3924 385 3976 394
rect 3976 385 3978 394
rect 4080 -295 4082 295
rect 4082 -295 4134 295
rect 4134 -295 4136 295
rect 4238 -394 4240 -385
rect 4240 -394 4292 -385
rect 4292 -394 4294 -385
rect 4238 -691 4294 -394
rect 4396 -295 4398 295
rect 4398 -295 4450 295
rect 4450 -295 4452 295
rect 4712 -295 4714 295
rect 4714 -295 4766 295
rect 4766 -295 4768 295
rect 4870 394 4926 691
rect 4870 385 4872 394
rect 4872 385 4924 394
rect 4924 385 4926 394
rect 5028 -295 5030 295
rect 5030 -295 5082 295
rect 5082 -295 5084 295
rect 5186 -394 5188 -385
rect 5188 -394 5240 -385
rect 5240 -394 5242 -385
rect 5186 -691 5242 -394
rect 5344 -295 5346 295
rect 5346 -295 5398 295
rect 5398 -295 5400 295
rect 5502 394 5558 691
rect 5502 385 5504 394
rect 5504 385 5556 394
rect 5556 385 5558 394
rect 5660 -295 5662 295
rect 5662 -295 5714 295
rect 5714 -295 5716 295
rect 5818 -394 5820 -385
rect 5820 -394 5872 -385
rect 5872 -394 5874 -385
rect 5818 -691 5874 -394
rect 5976 -295 5978 295
rect 5978 -295 6030 295
rect 6030 -295 6032 295
rect 6134 394 6190 691
rect 6134 385 6136 394
rect 6136 385 6188 394
rect 6188 385 6190 394
rect 6292 -295 6294 295
rect 6294 -295 6346 295
rect 6346 -295 6348 295
rect 6450 -394 6452 -385
rect 6452 -394 6504 -385
rect 6504 -394 6506 -385
rect 6450 -691 6506 -394
rect 6608 -295 6610 295
rect 6610 -295 6662 295
rect 6662 -295 6664 295
rect 6766 394 6822 691
rect 6766 385 6768 394
rect 6768 385 6820 394
rect 6820 385 6822 394
rect 6924 -295 6926 295
rect 6926 -295 6978 295
rect 6978 -295 6980 295
rect 7082 -394 7084 -385
rect 7084 -394 7136 -385
rect 7136 -394 7138 -385
rect 7082 -691 7138 -394
rect 7240 -295 7242 295
rect 7242 -295 7294 295
rect 7294 -295 7296 295
rect 7398 394 7454 691
rect 7398 385 7400 394
rect 7400 385 7452 394
rect 7452 385 7454 394
rect 7556 -295 7558 295
rect 7558 -295 7610 295
rect 7610 -295 7612 295
rect 7714 -394 7716 -385
rect 7716 -394 7768 -385
rect 7768 -394 7770 -385
rect 7714 -691 7770 -394
rect 7872 -295 7874 295
rect 7874 -295 7926 295
rect 7926 -295 7928 295
rect 8030 394 8086 691
rect 8030 385 8032 394
rect 8032 385 8084 394
rect 8084 385 8086 394
rect 8188 -295 8190 295
rect 8190 -295 8242 295
rect 8242 -295 8244 295
rect 8346 -394 8348 -385
rect 8348 -394 8400 -385
rect 8400 -394 8402 -385
rect 8346 -691 8402 -394
rect 8504 -295 8506 295
rect 8506 -295 8558 295
rect 8558 -295 8560 295
rect 8662 394 8718 691
rect 8662 385 8664 394
rect 8664 385 8716 394
rect 8716 385 8718 394
rect 8820 -295 8822 295
rect 8822 -295 8874 295
rect 8874 -295 8876 295
rect 8978 -394 8980 -385
rect 8980 -394 9032 -385
rect 9032 -394 9034 -385
rect 8978 -691 9034 -394
rect 9136 -295 9138 295
rect 9138 -295 9190 295
rect 9190 -295 9192 295
rect 9294 394 9350 691
rect 9294 385 9296 394
rect 9296 385 9348 394
rect 9348 385 9350 394
rect 9452 -295 9454 295
rect 9454 -295 9506 295
rect 9506 -295 9508 295
rect 9610 -394 9612 -385
rect 9612 -394 9664 -385
rect 9664 -394 9666 -385
rect 9610 -691 9666 -394
rect 9768 -295 9770 295
rect 9770 -295 9822 295
rect 9822 -295 9824 295
rect 9926 394 9982 691
rect 9926 385 9928 394
rect 9928 385 9980 394
rect 9980 385 9982 394
rect 10084 -295 10086 295
rect 10086 -295 10138 295
rect 10138 -295 10140 295
rect 10242 -394 10244 -385
rect 10244 -394 10296 -385
rect 10296 -394 10298 -385
rect 10242 -691 10298 -394
rect 10400 -295 10402 295
rect 10402 -295 10454 295
rect 10454 -295 10456 295
rect 10558 394 10614 691
rect 10558 385 10560 394
rect 10560 385 10612 394
rect 10612 385 10614 394
rect 10716 -295 10718 295
rect 10718 -295 10770 295
rect 10770 -295 10772 295
rect 10874 -394 10876 -385
rect 10876 -394 10928 -385
rect 10928 -394 10930 -385
rect 10874 -691 10930 -394
rect 11032 -295 11034 295
rect 11034 -295 11086 295
rect 11086 -295 11088 295
rect 11190 394 11246 691
rect 11190 385 11192 394
rect 11192 385 11244 394
rect 11244 385 11246 394
rect 11348 -295 11350 295
rect 11350 -295 11402 295
rect 11402 -295 11404 295
rect 11506 -394 11508 -385
rect 11508 -394 11560 -385
rect 11560 -394 11562 -385
rect 11506 -691 11562 -394
rect 11664 -295 11666 295
rect 11666 -295 11718 295
rect 11718 -295 11720 295
rect 11822 394 11878 691
rect 11822 385 11824 394
rect 11824 385 11876 394
rect 11876 385 11878 394
rect 11980 -295 11982 295
rect 11982 -295 12034 295
rect 12034 -295 12036 295
rect 12138 -394 12140 -385
rect 12140 -394 12192 -385
rect 12192 -394 12194 -385
rect 12138 -691 12194 -394
rect 12296 -295 12298 295
rect 12298 -295 12350 295
rect 12350 -295 12352 295
rect 12454 394 12510 691
rect 12454 385 12456 394
rect 12456 385 12508 394
rect 12508 385 12510 394
rect 12612 -295 12614 295
rect 12614 -295 12666 295
rect 12666 -295 12668 295
rect 12770 -394 12772 -385
rect 12772 -394 12824 -385
rect 12824 -394 12826 -385
rect 12770 -691 12826 -394
rect 12928 -295 12930 295
rect 12930 -295 12982 295
rect 12982 -295 12984 295
<< metal3 >>
rect -12989 691 12989 700
rect -12989 385 -12510 691
rect -12454 385 -11878 691
rect -11822 385 -11246 691
rect -11190 385 -10614 691
rect -10558 385 -9982 691
rect -9926 385 -9350 691
rect -9294 385 -8718 691
rect -8662 385 -8086 691
rect -8030 385 -7454 691
rect -7398 385 -6822 691
rect -6766 385 -6190 691
rect -6134 385 -5558 691
rect -5502 385 -4926 691
rect -4870 385 -3978 691
rect -3922 385 -3346 691
rect -3290 385 -2714 691
rect -2658 385 -2082 691
rect -2026 385 -1450 691
rect -1394 385 -818 691
rect -762 385 -186 691
rect -130 385 130 691
rect 186 385 762 691
rect 818 385 1394 691
rect 1450 385 2026 691
rect 2082 385 2658 691
rect 2714 385 3290 691
rect 3346 385 3922 691
rect 3978 385 4870 691
rect 4926 385 5502 691
rect 5558 385 6134 691
rect 6190 385 6766 691
rect 6822 385 7398 691
rect 7454 385 8030 691
rect 8086 385 8662 691
rect 8718 385 9294 691
rect 9350 385 9926 691
rect 9982 385 10558 691
rect 10614 385 11190 691
rect 11246 385 11822 691
rect 11878 385 12454 691
rect 12510 385 12989 691
rect -12989 380 12989 385
rect -12989 295 12989 300
rect -12989 -295 -12984 295
rect -12928 -295 -12668 295
rect -12612 -295 -12352 295
rect -12296 -295 -12036 295
rect -11980 -295 -11720 295
rect -11664 -295 -11404 295
rect -11348 -295 -11088 295
rect -11032 -295 -10772 295
rect -10716 -295 -10456 295
rect -10400 -295 -10140 295
rect -10084 -295 -9824 295
rect -9768 -295 -9508 295
rect -9452 -295 -9192 295
rect -9136 -295 -8876 295
rect -8820 -295 -8560 295
rect -8504 -295 -8244 295
rect -8188 -295 -7928 295
rect -7872 -295 -7612 295
rect -7556 -295 -7296 295
rect -7240 -295 -6980 295
rect -6924 -295 -6664 295
rect -6608 -295 -6348 295
rect -6292 -295 -6032 295
rect -5976 -295 -5716 295
rect -5660 -295 -5400 295
rect -5344 -295 -5084 295
rect -5028 -295 -4768 295
rect -4712 -295 -4452 295
rect -4396 -295 -4136 295
rect -4080 -295 -3820 295
rect -3764 -295 -3504 295
rect -3448 -295 -3188 295
rect -3132 -295 -2872 295
rect -2816 -295 -2556 295
rect -2500 -295 -2240 295
rect -2184 -295 -1924 295
rect -1868 -295 -1608 295
rect -1552 -295 -1292 295
rect -1236 -295 -976 295
rect -920 -295 -660 295
rect -604 -295 -344 295
rect -288 -295 -28 295
rect 28 -295 288 295
rect 344 -295 604 295
rect 660 -295 920 295
rect 976 -295 1236 295
rect 1292 -295 1552 295
rect 1608 -295 1868 295
rect 1924 -295 2184 295
rect 2240 -295 2500 295
rect 2556 -295 2816 295
rect 2872 -295 3132 295
rect 3188 -295 3448 295
rect 3504 -295 3764 295
rect 3820 -295 4080 295
rect 4136 -295 4396 295
rect 4452 -295 4712 295
rect 4768 -295 5028 295
rect 5084 -295 5344 295
rect 5400 -295 5660 295
rect 5716 -295 5976 295
rect 6032 -295 6292 295
rect 6348 -295 6608 295
rect 6664 -295 6924 295
rect 6980 -295 7240 295
rect 7296 -295 7556 295
rect 7612 -295 7872 295
rect 7928 -295 8188 295
rect 8244 -295 8504 295
rect 8560 -295 8820 295
rect 8876 -295 9136 295
rect 9192 -295 9452 295
rect 9508 -295 9768 295
rect 9824 -295 10084 295
rect 10140 -295 10400 295
rect 10456 -295 10716 295
rect 10772 -295 11032 295
rect 11088 -295 11348 295
rect 11404 -295 11664 295
rect 11720 -295 11980 295
rect 12036 -295 12296 295
rect 12352 -295 12612 295
rect 12668 -295 12928 295
rect 12984 -295 12989 295
rect -12989 -300 12989 -295
rect -12989 -385 12989 -380
rect -12989 -691 -12826 -385
rect -12770 -691 -12194 -385
rect -12138 -691 -11562 -385
rect -11506 -691 -10930 -385
rect -10874 -691 -10298 -385
rect -10242 -691 -9666 -385
rect -9610 -691 -9034 -385
rect -8978 -691 -8402 -385
rect -8346 -691 -7770 -385
rect -7714 -691 -7138 -385
rect -7082 -691 -6506 -385
rect -6450 -691 -5874 -385
rect -5818 -691 -5242 -385
rect -5186 -691 -4294 -385
rect -4238 -691 -3662 -385
rect -3606 -691 -3030 -385
rect -2974 -691 -2398 -385
rect -2342 -691 -1766 -385
rect -1710 -691 -1134 -385
rect -1078 -691 -502 -385
rect -446 -691 446 -385
rect 502 -691 1078 -385
rect 1134 -691 1710 -385
rect 1766 -691 2342 -385
rect 2398 -691 2974 -385
rect 3030 -691 3606 -385
rect 3662 -691 4238 -385
rect 4294 -691 5186 -385
rect 5242 -691 5818 -385
rect 5874 -691 6450 -385
rect 6506 -691 7082 -385
rect 7138 -691 7714 -385
rect 7770 -691 8346 -385
rect 8402 -691 8978 -385
rect 9034 -691 9610 -385
rect 9666 -691 10242 -385
rect 10298 -691 10874 -385
rect 10930 -691 11506 -385
rect 11562 -691 12138 -385
rect 12194 -691 12770 -385
rect 12826 -691 12989 -385
rect -12989 -700 12989 -691
<< properties >>
string FIXED_BBOX -13090 -393 13090 393
string gencell sky130_fd_pr__nfet_g5v0d10v5
string library sky130
string parameters w 2 l 0.5 m 1 nf 164 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
